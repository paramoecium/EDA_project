module top ( PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D );
input PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D;
wire n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241;
buf ( n243 , n2315 );
buf ( n244 , n2317 );
buf ( n245 , n2319 );
buf ( n246 , n2321 );
buf ( n247 , n2323 );
buf ( n248 , n2325 );
buf ( n249 , n2327 );
buf ( n250 , n2329 );
buf ( n251 , n2331 );
buf ( n252 , n2333 );
buf ( n253 , n2335 );
buf ( n254 , n2337 );
buf ( n255 , n2339 );
buf ( n256 , n2341 );
buf ( n257 , n2343 );
buf ( n258 , n2345 );
buf ( n259 , n2347 );
buf ( n260 , n2349 );
buf ( n261 , n2351 );
buf ( n262 , n2353 );
buf ( n263 , n2355 );
buf ( n264 , n2357 );
buf ( n265 , n2359 );
buf ( n266 , n2361 );
buf ( n267 , n2363 );
buf ( n268 , n2365 );
buf ( n269 , n2367 );
buf ( n270 , n2369 );
buf ( n271 , n2371 );
buf ( n272 , n2373 );
buf ( n273 , n2375 );
buf ( n274 , n2377 );
buf ( n275 , n2379 );
buf ( n276 , n2381 );
buf ( n277 , n2383 );
buf ( n278 , n2385 );
buf ( n279 , n2387 );
buf ( n280 , n2389 );
buf ( n281 , n2391 );
buf ( n282 , n2393 );
buf ( n283 , n2395 );
buf ( n284 , n2397 );
buf ( n285 , n2399 );
buf ( n286 , n2401 );
buf ( n287 , n2403 );
buf ( n288 , n2405 );
buf ( n289 , n2407 );
buf ( n290 , n2409 );
buf ( n291 , n2411 );
buf ( n292 , n2413 );
buf ( n293 , n2415 );
buf ( n294 , n2417 );
buf ( PO_rd , n2419 );
buf ( PO_wr , n2421 );
buf ( DFF_state_reg_S , n2425 );
buf ( DFF_state_reg_R , n2426 );
buf ( DFF_state_reg_CK , n2427 );
buf ( DFF_state_reg_D , n2429 );
buf ( n295 , n2431 );
buf ( n296 , n2432 );
buf ( n297 , n2433 );
buf ( n298 , n2437 );
buf ( n299 , n2439 );
buf ( n300 , n2440 );
buf ( n301 , n2441 );
buf ( n302 , n2453 );
buf ( n303 , n2455 );
buf ( n304 , n2456 );
buf ( n305 , n2457 );
buf ( n306 , n2468 );
buf ( n307 , n2470 );
buf ( n308 , n2471 );
buf ( n309 , n2472 );
buf ( n310 , n2483 );
buf ( n311 , n2485 );
buf ( n312 , n2486 );
buf ( n313 , n2487 );
buf ( n314 , n2498 );
buf ( n315 , n2500 );
buf ( n316 , n2501 );
buf ( n317 , n2502 );
buf ( n318 , n2513 );
buf ( n319 , n2515 );
buf ( n320 , n2516 );
buf ( n321 , n2517 );
buf ( n322 , n2528 );
buf ( n323 , n2530 );
buf ( n324 , n2531 );
buf ( n325 , n2532 );
buf ( n326 , n2543 );
buf ( n327 , n2545 );
buf ( n328 , n2546 );
buf ( n329 , n2547 );
buf ( n330 , n2558 );
buf ( n331 , n2560 );
buf ( n332 , n2561 );
buf ( n333 , n2562 );
buf ( n334 , n2573 );
buf ( n335 , n2575 );
buf ( n336 , n2576 );
buf ( n337 , n2577 );
buf ( n338 , n2588 );
buf ( n339 , n2590 );
buf ( n340 , n2591 );
buf ( n341 , n2592 );
buf ( n342 , n2603 );
buf ( n343 , n2605 );
buf ( n344 , n2606 );
buf ( n345 , n2607 );
buf ( n346 , n2618 );
buf ( n347 , n2620 );
buf ( n348 , n2621 );
buf ( n349 , n2622 );
buf ( n350 , n2633 );
buf ( n351 , n2635 );
buf ( n352 , n2636 );
buf ( n353 , n2637 );
buf ( n354 , n2648 );
buf ( n355 , n2650 );
buf ( n356 , n2651 );
buf ( n357 , n2652 );
buf ( n358 , n2663 );
buf ( n359 , n2665 );
buf ( n360 , n2666 );
buf ( n361 , n2667 );
buf ( n362 , n2678 );
buf ( n363 , n2680 );
buf ( n364 , n2681 );
buf ( n365 , n2682 );
buf ( n366 , n2693 );
buf ( n367 , n2695 );
buf ( n368 , n2696 );
buf ( n369 , n2697 );
buf ( n370 , n2708 );
buf ( n371 , n2710 );
buf ( n372 , n2711 );
buf ( n373 , n2712 );
buf ( n374 , n2723 );
buf ( n375 , n2725 );
buf ( n376 , n2726 );
buf ( n377 , n2727 );
buf ( n378 , n2738 );
buf ( n379 , n2740 );
buf ( n380 , n2741 );
buf ( n381 , n2742 );
buf ( n382 , n2753 );
buf ( n383 , n2755 );
buf ( n384 , n2756 );
buf ( n385 , n2757 );
buf ( n386 , n2768 );
buf ( n387 , n2770 );
buf ( n388 , n2771 );
buf ( n389 , n2772 );
buf ( n390 , n2783 );
buf ( n391 , n2785 );
buf ( n392 , n2786 );
buf ( n393 , n2787 );
buf ( n394 , n2798 );
buf ( n395 , n2800 );
buf ( n396 , n2801 );
buf ( n397 , n2802 );
buf ( n398 , n2813 );
buf ( n399 , n2815 );
buf ( n400 , n2816 );
buf ( n401 , n2817 );
buf ( n402 , n2828 );
buf ( n403 , n2830 );
buf ( n404 , n2831 );
buf ( n405 , n2832 );
buf ( n406 , n2843 );
buf ( n407 , n2845 );
buf ( n408 , n2846 );
buf ( n409 , n2847 );
buf ( n410 , n2858 );
buf ( n411 , n2860 );
buf ( n412 , n2861 );
buf ( n413 , n2862 );
buf ( n414 , n2873 );
buf ( n415 , n2875 );
buf ( n416 , n2876 );
buf ( n417 , n2877 );
buf ( n418 , n2888 );
buf ( n419 , n2889 );
buf ( n420 , n2890 );
buf ( n421 , n2891 );
buf ( n422 , n2903 );
buf ( n423 , n2905 );
buf ( n424 , n2906 );
buf ( n425 , n2907 );
buf ( n426 , n3311 );
buf ( n427 , n3313 );
buf ( n428 , n3314 );
buf ( n429 , n3315 );
buf ( n430 , n3355 );
buf ( n431 , n3357 );
buf ( n432 , n3358 );
buf ( n433 , n3359 );
buf ( n434 , n6733 );
buf ( n435 , n6734 );
buf ( n436 , n6735 );
buf ( n437 , n6736 );
buf ( n438 , n7089 );
buf ( n439 , n7090 );
buf ( n440 , n7091 );
buf ( n441 , n7092 );
buf ( n442 , n7163 );
buf ( n443 , n7164 );
buf ( n444 , n7165 );
buf ( n445 , n7166 );
buf ( n446 , n7237 );
buf ( n447 , n7238 );
buf ( n448 , n7239 );
buf ( n449 , n7240 );
buf ( n450 , n7311 );
buf ( n451 , n7312 );
buf ( n452 , n7313 );
buf ( n453 , n7314 );
buf ( n454 , n7385 );
buf ( n455 , n7386 );
buf ( n456 , n7387 );
buf ( n457 , n7388 );
buf ( n458 , n7459 );
buf ( n459 , n7460 );
buf ( n460 , n7461 );
buf ( n461 , n7462 );
buf ( n462 , n7533 );
buf ( n463 , n7534 );
buf ( n464 , n7535 );
buf ( n465 , n7536 );
buf ( n466 , n7607 );
buf ( n467 , n7608 );
buf ( n468 , n7609 );
buf ( n469 , n7610 );
buf ( n470 , n7681 );
buf ( n471 , n7682 );
buf ( n472 , n7683 );
buf ( n473 , n7684 );
buf ( n474 , n7755 );
buf ( n475 , n7756 );
buf ( n476 , n7757 );
buf ( n477 , n7758 );
buf ( n478 , n7829 );
buf ( n479 , n7830 );
buf ( n480 , n7831 );
buf ( n481 , n7832 );
buf ( n482 , n7903 );
buf ( n483 , n7904 );
buf ( n484 , n7905 );
buf ( n485 , n7906 );
buf ( n486 , n7977 );
buf ( n487 , n7978 );
buf ( n488 , n7979 );
buf ( n489 , n7980 );
buf ( n490 , n8051 );
buf ( n491 , n8052 );
buf ( n492 , n8053 );
buf ( n493 , n8054 );
buf ( n494 , n8125 );
buf ( n495 , n8126 );
buf ( n496 , n8127 );
buf ( n497 , n8128 );
buf ( n498 , n8199 );
buf ( n499 , n8200 );
buf ( n500 , n8201 );
buf ( n501 , n8202 );
buf ( n502 , n8273 );
buf ( n503 , n8274 );
buf ( n504 , n8275 );
buf ( n505 , n8276 );
buf ( n506 , n8347 );
buf ( n507 , n8348 );
buf ( n508 , n8349 );
buf ( n509 , n8350 );
buf ( n510 , n8421 );
buf ( n511 , n8422 );
buf ( n512 , n8423 );
buf ( n513 , n8424 );
buf ( n514 , n8495 );
buf ( n515 , n8496 );
buf ( n516 , n8497 );
buf ( n517 , n8498 );
buf ( n518 , n8569 );
buf ( n519 , n8570 );
buf ( n520 , n8571 );
buf ( n521 , n8572 );
buf ( n522 , n8643 );
buf ( n523 , n8644 );
buf ( n524 , n8645 );
buf ( n525 , n8646 );
buf ( n526 , n8717 );
buf ( n527 , n8718 );
buf ( n528 , n8719 );
buf ( n529 , n8720 );
buf ( n530 , n8791 );
buf ( n531 , n8792 );
buf ( n532 , n8793 );
buf ( n533 , n8794 );
buf ( n534 , n8865 );
buf ( n535 , n8866 );
buf ( n536 , n8867 );
buf ( n537 , n8868 );
buf ( n538 , n8939 );
buf ( n539 , n8940 );
buf ( n540 , n8941 );
buf ( n541 , n8942 );
buf ( n542 , n9013 );
buf ( n543 , n9014 );
buf ( n544 , n9015 );
buf ( n545 , n9016 );
buf ( n546 , n9087 );
buf ( n547 , n9088 );
buf ( n548 , n9089 );
buf ( n549 , n9090 );
buf ( n550 , n9124 );
buf ( n551 , n9125 );
buf ( n552 , n9126 );
buf ( n553 , n9127 );
buf ( n554 , n9157 );
buf ( n555 , n9158 );
buf ( n556 , n9159 );
buf ( n557 , n9160 );
buf ( n558 , n9190 );
buf ( n559 , n9191 );
buf ( n560 , n9192 );
buf ( n561 , n9193 );
buf ( n562 , n9223 );
buf ( n563 , n9224 );
buf ( n564 , n9225 );
buf ( n565 , n9226 );
buf ( n566 , n9256 );
buf ( n567 , n9257 );
buf ( n568 , n9258 );
buf ( n569 , n9259 );
buf ( n570 , n9289 );
buf ( n571 , n9290 );
buf ( n572 , n9291 );
buf ( n573 , n9292 );
buf ( n574 , n9322 );
buf ( n575 , n9323 );
buf ( n576 , n9324 );
buf ( n577 , n9325 );
buf ( n578 , n9355 );
buf ( n579 , n9356 );
buf ( n580 , n9357 );
buf ( n581 , n9358 );
buf ( n582 , n9388 );
buf ( n583 , n9389 );
buf ( n584 , n9390 );
buf ( n585 , n9391 );
buf ( n586 , n9421 );
buf ( n587 , n9422 );
buf ( n588 , n9423 );
buf ( n589 , n9424 );
buf ( n590 , n9454 );
buf ( n591 , n9455 );
buf ( n592 , n9456 );
buf ( n593 , n9457 );
buf ( n594 , n9487 );
buf ( n595 , n9488 );
buf ( n596 , n9489 );
buf ( n597 , n9490 );
buf ( n598 , n9520 );
buf ( n599 , n9521 );
buf ( n600 , n9522 );
buf ( n601 , n9523 );
buf ( n602 , n9553 );
buf ( n603 , n9554 );
buf ( n604 , n9555 );
buf ( n605 , n9556 );
buf ( n606 , n9586 );
buf ( n607 , n9587 );
buf ( n608 , n9588 );
buf ( n609 , n9589 );
buf ( n610 , n9619 );
buf ( n611 , n9620 );
buf ( n612 , n9621 );
buf ( n613 , n9622 );
buf ( n614 , n9652 );
buf ( n615 , n9653 );
buf ( n616 , n9654 );
buf ( n617 , n9655 );
buf ( n618 , n9685 );
buf ( n619 , n9686 );
buf ( n620 , n9687 );
buf ( n621 , n9688 );
buf ( n622 , n9718 );
buf ( n623 , n9719 );
buf ( n624 , n9720 );
buf ( n625 , n9721 );
buf ( n626 , n9751 );
buf ( n627 , n9752 );
buf ( n628 , n9753 );
buf ( n629 , n9754 );
buf ( n630 , n9784 );
buf ( n631 , n9785 );
buf ( n632 , n9786 );
buf ( n633 , n9787 );
buf ( n634 , n9817 );
buf ( n635 , n9818 );
buf ( n636 , n9819 );
buf ( n637 , n9820 );
buf ( n638 , n9850 );
buf ( n639 , n9851 );
buf ( n640 , n9852 );
buf ( n641 , n9853 );
buf ( n642 , n9883 );
buf ( n643 , n9884 );
buf ( n644 , n9885 );
buf ( n645 , n9886 );
buf ( n646 , n9916 );
buf ( n647 , n9917 );
buf ( n648 , n9918 );
buf ( n649 , n9919 );
buf ( n650 , n9949 );
buf ( n651 , n9950 );
buf ( n652 , n9951 );
buf ( n653 , n9952 );
buf ( n654 , n9982 );
buf ( n655 , n9983 );
buf ( n656 , n9984 );
buf ( n657 , n9985 );
buf ( n658 , n10015 );
buf ( n659 , n10016 );
buf ( n660 , n10017 );
buf ( n661 , n10018 );
buf ( n662 , n10048 );
buf ( n663 , n10049 );
buf ( n664 , n10050 );
buf ( n665 , n10051 );
buf ( n666 , n10124 );
buf ( n667 , n10125 );
buf ( n668 , n10126 );
buf ( n669 , n10127 );
buf ( n670 , n10189 );
buf ( n671 , n10190 );
buf ( n672 , n10191 );
buf ( n673 , n10192 );
buf ( n674 , n10229 );
buf ( n675 , n10230 );
buf ( n676 , n10231 );
buf ( n677 , n10232 );
buf ( n678 , n10265 );
buf ( n679 , n10266 );
buf ( n680 , n10267 );
buf ( n681 , n10268 );
buf ( n682 , n10298 );
buf ( n683 , n10299 );
buf ( n684 , n10300 );
buf ( n685 , n10301 );
buf ( n686 , n10331 );
buf ( n687 , n10332 );
buf ( n688 , n10333 );
buf ( n689 , n10334 );
buf ( n690 , n10364 );
buf ( n691 , n10365 );
buf ( n692 , n10366 );
buf ( n693 , n10367 );
buf ( n694 , n10397 );
buf ( n695 , n10398 );
buf ( n696 , n10399 );
buf ( n697 , n10400 );
buf ( n698 , n10430 );
buf ( n699 , n10431 );
buf ( n700 , n10432 );
buf ( n701 , n10433 );
buf ( n702 , n10463 );
buf ( n703 , n10464 );
buf ( n704 , n10465 );
buf ( n705 , n10466 );
buf ( n706 , n10496 );
buf ( n707 , n10497 );
buf ( n708 , n10498 );
buf ( n709 , n10499 );
buf ( n710 , n10529 );
buf ( n711 , n10530 );
buf ( n712 , n10531 );
buf ( n713 , n10532 );
buf ( n714 , n10562 );
buf ( n715 , n10563 );
buf ( n716 , n10564 );
buf ( n717 , n10565 );
buf ( n718 , n10595 );
buf ( n719 , n10596 );
buf ( n720 , n10597 );
buf ( n721 , n10598 );
buf ( n722 , n10628 );
buf ( n723 , n10629 );
buf ( n724 , n10630 );
buf ( n725 , n10631 );
buf ( n726 , n10661 );
buf ( n727 , n10662 );
buf ( n728 , n10663 );
buf ( n729 , n10664 );
buf ( n730 , n10694 );
buf ( n731 , n10695 );
buf ( n732 , n10696 );
buf ( n733 , n10697 );
buf ( n734 , n10727 );
buf ( n735 , n10728 );
buf ( n736 , n10729 );
buf ( n737 , n10730 );
buf ( n738 , n10760 );
buf ( n739 , n10761 );
buf ( n740 , n10762 );
buf ( n741 , n10763 );
buf ( n742 , n10793 );
buf ( n743 , n10794 );
buf ( n744 , n10795 );
buf ( n745 , n10796 );
buf ( n746 , n10826 );
buf ( n747 , n10827 );
buf ( n748 , n10828 );
buf ( n749 , n10829 );
buf ( n750 , n10859 );
buf ( n751 , n10860 );
buf ( n752 , n10861 );
buf ( n753 , n10862 );
buf ( n754 , n10892 );
buf ( n755 , n10893 );
buf ( n756 , n10894 );
buf ( n757 , n10895 );
buf ( n758 , n10925 );
buf ( n759 , n10926 );
buf ( n760 , n10927 );
buf ( n761 , n10928 );
buf ( n762 , n10958 );
buf ( n763 , n10959 );
buf ( n764 , n10960 );
buf ( n765 , n10961 );
buf ( n766 , n10991 );
buf ( n767 , n10992 );
buf ( n768 , n10993 );
buf ( n769 , n10994 );
buf ( n770 , n11024 );
buf ( n771 , n11025 );
buf ( n772 , n11026 );
buf ( n773 , n11027 );
buf ( n774 , n11057 );
buf ( n775 , n11058 );
buf ( n776 , n11059 );
buf ( n777 , n11060 );
buf ( n778 , n11090 );
buf ( n779 , n11091 );
buf ( n780 , n11092 );
buf ( n781 , n11093 );
buf ( n782 , n11123 );
buf ( n783 , n11124 );
buf ( n784 , n11125 );
buf ( n785 , n11126 );
buf ( n786 , n11156 );
buf ( n787 , n11157 );
buf ( n788 , n11158 );
buf ( n789 , n11159 );
buf ( n790 , n11189 );
buf ( n791 , n11190 );
buf ( n792 , n11191 );
buf ( n793 , n11192 );
buf ( n794 , n11222 );
buf ( n795 , n11223 );
buf ( n796 , n11224 );
buf ( n797 , n11225 );
buf ( n798 , n11255 );
buf ( n799 , n11256 );
buf ( n800 , n11257 );
buf ( n801 , n11258 );
buf ( n802 , n11284 );
buf ( DFF_B_reg_S , n11285 );
buf ( DFF_B_reg_R , n11286 );
buf ( DFF_B_reg_CK , n11287 );
buf ( DFF_B_reg_D , n11901 );
buf ( n803 , n11902 );
buf ( n804 , n11903 );
buf ( n805 , n11904 );
buf ( n806 , n11937 );
buf ( n807 , n11938 );
buf ( n808 , n11939 );
buf ( n809 , n11940 );
buf ( n810 , n11971 );
buf ( n811 , n11972 );
buf ( n812 , n11973 );
buf ( n813 , n11974 );
buf ( n814 , n12005 );
buf ( n815 , n12006 );
buf ( n816 , n12007 );
buf ( n817 , n12008 );
buf ( n818 , n12039 );
buf ( n819 , n12040 );
buf ( n820 , n12041 );
buf ( n821 , n12042 );
buf ( n822 , n12073 );
buf ( n823 , n12074 );
buf ( n824 , n12075 );
buf ( n825 , n12076 );
buf ( n826 , n12107 );
buf ( n827 , n12108 );
buf ( n828 , n12109 );
buf ( n829 , n12110 );
buf ( n830 , n12141 );
buf ( n831 , n12142 );
buf ( n832 , n12143 );
buf ( n833 , n12144 );
buf ( n834 , n12175 );
buf ( n835 , n12176 );
buf ( n836 , n12177 );
buf ( n837 , n12178 );
buf ( n838 , n12209 );
buf ( n839 , n12210 );
buf ( n840 , n12211 );
buf ( n841 , n12212 );
buf ( n842 , n12243 );
buf ( n843 , n12244 );
buf ( n844 , n12245 );
buf ( n845 , n12246 );
buf ( n846 , n12277 );
buf ( n847 , n12278 );
buf ( n848 , n12279 );
buf ( n849 , n12280 );
buf ( n850 , n12311 );
buf ( n851 , n12312 );
buf ( n852 , n12313 );
buf ( n853 , n12314 );
buf ( n854 , n12345 );
buf ( n855 , n12346 );
buf ( n856 , n12347 );
buf ( n857 , n12348 );
buf ( n858 , n12379 );
buf ( n859 , n12380 );
buf ( n860 , n12381 );
buf ( n861 , n12382 );
buf ( n862 , n12413 );
buf ( n863 , n12414 );
buf ( n864 , n12415 );
buf ( n865 , n12416 );
buf ( n866 , n12447 );
buf ( n867 , n12448 );
buf ( n868 , n12449 );
buf ( n869 , n12450 );
buf ( n870 , n12481 );
buf ( n871 , n12482 );
buf ( n872 , n12483 );
buf ( n873 , n12484 );
buf ( n874 , n12515 );
buf ( n875 , n12516 );
buf ( n876 , n12517 );
buf ( n877 , n12518 );
buf ( n878 , n12549 );
buf ( n879 , n12550 );
buf ( n880 , n12551 );
buf ( n881 , n12552 );
buf ( n882 , n12583 );
buf ( n883 , n12584 );
buf ( n884 , n12585 );
buf ( n885 , n12586 );
buf ( n886 , n12617 );
buf ( n887 , n12618 );
buf ( n888 , n12619 );
buf ( n889 , n12620 );
buf ( n890 , n12651 );
buf ( n891 , n12652 );
buf ( n892 , n12653 );
buf ( n893 , n12654 );
buf ( n894 , n12685 );
buf ( n895 , n12686 );
buf ( n896 , n12687 );
buf ( n897 , n12688 );
buf ( n898 , n12719 );
buf ( n899 , n12720 );
buf ( n900 , n12721 );
buf ( n901 , n12722 );
buf ( n902 , n12753 );
buf ( n903 , n12754 );
buf ( n904 , n12755 );
buf ( n905 , n12756 );
buf ( n906 , n12787 );
buf ( n907 , n12788 );
buf ( n908 , n12789 );
buf ( n909 , n12790 );
buf ( n910 , n12821 );
buf ( n911 , n12822 );
buf ( n912 , n12823 );
buf ( n913 , n12824 );
buf ( n914 , n12855 );
buf ( n915 , n12856 );
buf ( n916 , n12857 );
buf ( n917 , n12858 );
buf ( n918 , n12889 );
buf ( n919 , n12890 );
buf ( n920 , n12891 );
buf ( n921 , n12892 );
buf ( n922 , n12923 );
buf ( n923 , n12924 );
buf ( n924 , n12925 );
buf ( n925 , n12926 );
buf ( n926 , n12956 );
buf ( n927 , n12957 );
buf ( n928 , n12958 );
buf ( n929 , n12959 );
buf ( n930 , n12985 );
buf ( n931 , n12986 );
buf ( n932 , n12987 );
buf ( n933 , n12988 );
buf ( n934 , n13677 );
buf ( n935 , n13678 );
buf ( n936 , n13679 );
buf ( n937 , n13680 );
buf ( n938 , n13718 );
buf ( n939 , n13719 );
buf ( n940 , n13720 );
buf ( n941 , n13721 );
buf ( n942 , n14169 );
buf ( n943 , n14170 );
buf ( n944 , n14171 );
buf ( n945 , n14172 );
buf ( n946 , n14210 );
buf ( n947 , n14211 );
buf ( n948 , n14212 );
buf ( n949 , n14213 );
buf ( n950 , n14252 );
buf ( n951 , n14253 );
buf ( n952 , n14254 );
buf ( n953 , n14255 );
buf ( n954 , n14293 );
buf ( n955 , n14294 );
buf ( n956 , n14295 );
buf ( n957 , n14296 );
buf ( n958 , n14334 );
buf ( n959 , n14335 );
buf ( n960 , n14336 );
buf ( n961 , n14337 );
buf ( n962 , n14375 );
buf ( n963 , n14376 );
buf ( n964 , n14377 );
buf ( n965 , n14378 );
buf ( n966 , n14416 );
buf ( n967 , n14417 );
buf ( n968 , n14418 );
buf ( n969 , n14419 );
buf ( n970 , n14457 );
buf ( n971 , n14458 );
buf ( n972 , n14459 );
buf ( n973 , n14460 );
buf ( n974 , n14498 );
buf ( n975 , n14499 );
buf ( n976 , n14500 );
buf ( n977 , n14501 );
buf ( n978 , n14539 );
buf ( n979 , n14540 );
buf ( n980 , n14541 );
buf ( n981 , n14542 );
buf ( n982 , n14580 );
buf ( n983 , n14581 );
buf ( n984 , n14582 );
buf ( n985 , n14583 );
buf ( n986 , n14621 );
buf ( n987 , n14622 );
buf ( n988 , n14623 );
buf ( n989 , n14624 );
buf ( n990 , n14662 );
buf ( n991 , n14663 );
buf ( n992 , n14664 );
buf ( n993 , n14665 );
buf ( n994 , n14703 );
buf ( n995 , n14704 );
buf ( n996 , n14705 );
buf ( n997 , n14706 );
buf ( n998 , n14744 );
buf ( n999 , n14745 );
buf ( n1000 , n14746 );
buf ( n1001 , n14747 );
buf ( n1002 , n14785 );
buf ( n1003 , n14786 );
buf ( n1004 , n14787 );
buf ( n1005 , n14788 );
buf ( n1006 , n14826 );
buf ( n1007 , n14827 );
buf ( n1008 , n14828 );
buf ( n1009 , n14829 );
buf ( n1010 , n14867 );
buf ( n1011 , n14868 );
buf ( n1012 , n14869 );
buf ( n1013 , n14870 );
buf ( n1014 , n14880 );
buf ( n1015 , n14881 );
buf ( n1016 , n14882 );
buf ( n1017 , n14883 );
buf ( n1018 , n14891 );
buf ( n1019 , n14892 );
buf ( n1020 , n14893 );
buf ( n1021 , n14894 );
buf ( n1022 , n14902 );
buf ( n1023 , n14903 );
buf ( n1024 , n14904 );
buf ( n1025 , n14905 );
buf ( n1026 , n14913 );
buf ( n1027 , n14914 );
buf ( n1028 , n14915 );
buf ( n1029 , n14916 );
buf ( n1030 , n14924 );
buf ( n1031 , n14925 );
buf ( n1032 , n14926 );
buf ( n1033 , n14927 );
buf ( n1034 , n14935 );
buf ( n1035 , n14936 );
buf ( n1036 , n14937 );
buf ( n1037 , n14938 );
buf ( n1038 , n14946 );
buf ( n1039 , n14947 );
buf ( n1040 , n14948 );
buf ( n1041 , n14949 );
buf ( n1042 , n14957 );
buf ( n1043 , n14958 );
buf ( n1044 , n14959 );
buf ( n1045 , n14960 );
buf ( n1046 , n14968 );
buf ( n1047 , n14969 );
buf ( n1048 , n14970 );
buf ( n1049 , n14971 );
buf ( n1050 , n14979 );
buf ( n1051 , n14980 );
buf ( n1052 , n14981 );
buf ( n1053 , n14982 );
buf ( n1054 , n14990 );
buf ( n1055 , n14991 );
buf ( n1056 , n14992 );
buf ( n1057 , n14993 );
buf ( n1058 , n15001 );
buf ( n1059 , n15002 );
buf ( n1060 , n15003 );
buf ( n1061 , n15004 );
buf ( n1062 , n15012 );
buf ( n1063 , n15013 );
buf ( n1064 , n15014 );
buf ( n1065 , n15015 );
buf ( n1066 , n15023 );
buf ( n1067 , n15024 );
buf ( n1068 , n15025 );
buf ( n1069 , n15026 );
buf ( n1070 , n15034 );
buf ( n1071 , n15035 );
buf ( n1072 , n15036 );
buf ( n1073 , n15037 );
buf ( n1074 , n15045 );
buf ( n1075 , n15046 );
buf ( n1076 , n15047 );
buf ( n1077 , n15048 );
buf ( n1078 , n15056 );
buf ( n1079 , n15057 );
buf ( n1080 , n15058 );
buf ( n1081 , n15059 );
buf ( n1082 , n15067 );
buf ( n1083 , n15068 );
buf ( n1084 , n15069 );
buf ( n1085 , n15070 );
buf ( n1086 , n15078 );
buf ( n1087 , n15079 );
buf ( n1088 , n15080 );
buf ( n1089 , n15081 );
buf ( n1090 , n15089 );
buf ( n1091 , n15090 );
buf ( n1092 , n15091 );
buf ( n1093 , n15092 );
buf ( n1094 , n15100 );
buf ( n1095 , n15101 );
buf ( n1096 , n15102 );
buf ( n1097 , n15103 );
buf ( n1098 , n15111 );
buf ( n1099 , n15112 );
buf ( n1100 , n15113 );
buf ( n1101 , n15114 );
buf ( n1102 , n15122 );
buf ( n1103 , n15123 );
buf ( n1104 , n15124 );
buf ( n1105 , n15125 );
buf ( n1106 , n15133 );
buf ( n1107 , n15134 );
buf ( n1108 , n15135 );
buf ( n1109 , n15136 );
buf ( n1110 , n15144 );
buf ( n1111 , n15145 );
buf ( n1112 , n15146 );
buf ( n1113 , n15147 );
buf ( n1114 , n15155 );
buf ( n1115 , n15156 );
buf ( n1116 , n15157 );
buf ( n1117 , n15158 );
buf ( n1118 , n15166 );
buf ( n1119 , n15167 );
buf ( n1120 , n15168 );
buf ( n1121 , n15169 );
buf ( n1122 , n15177 );
buf ( n1123 , n15178 );
buf ( n1124 , n15179 );
buf ( n1125 , n15180 );
buf ( n1126 , n15188 );
buf ( n1127 , n15189 );
buf ( n1128 , n15190 );
buf ( n1129 , n15191 );
buf ( n1130 , n15199 );
buf ( n1131 , n15200 );
buf ( n1132 , n15201 );
buf ( n1133 , n15202 );
buf ( n1134 , n15210 );
buf ( n1135 , n15211 );
buf ( n1136 , n15212 );
buf ( n1137 , n15213 );
buf ( n1138 , n15221 );
buf ( DFF_rd_reg_S , n15222 );
buf ( DFF_rd_reg_R , n15223 );
buf ( DFF_rd_reg_CK , n15224 );
buf ( DFF_rd_reg_D , n15234 );
buf ( DFF_wr_reg_S , n15235 );
buf ( DFF_wr_reg_R , n15236 );
buf ( DFF_wr_reg_CK , n15237 );
buf ( DFF_wr_reg_D , n15241 );
buf ( n2280 , PI_clock );
buf ( n2281 , PI_reset );
buf ( n2282 , n0 );
buf ( n2283 , n1 );
buf ( n2284 , n2 );
buf ( n2285 , n3 );
buf ( n2286 , n4 );
buf ( n2287 , n5 );
buf ( n2288 , n6 );
buf ( n2289 , n7 );
buf ( n2290 , n8 );
buf ( n2291 , n9 );
buf ( n2292 , n10 );
buf ( n2293 , n11 );
buf ( n2294 , n12 );
buf ( n2295 , n13 );
buf ( n2296 , n14 );
buf ( n2297 , n15 );
buf ( n2298 , n16 );
buf ( n2299 , n17 );
buf ( n2300 , n18 );
buf ( n2301 , n19 );
buf ( n2302 , n20 );
buf ( n2303 , n21 );
buf ( n2304 , n22 );
buf ( n2305 , n23 );
buf ( n2306 , n24 );
buf ( n2307 , n25 );
buf ( n2308 , n26 );
buf ( n2309 , n27 );
buf ( n2310 , n28 );
buf ( n2311 , n29 );
buf ( n2312 , n30 );
buf ( n2313 , n31 );
buf ( n2314 , n210 );
buf ( n2315 , n2314 );
buf ( n2316 , n209 );
buf ( n2317 , n2316 );
buf ( n2318 , n208 );
buf ( n2319 , n2318 );
buf ( n2320 , n207 );
buf ( n2321 , n2320 );
buf ( n2322 , n206 );
buf ( n2323 , n2322 );
buf ( n2324 , n205 );
buf ( n2325 , n2324 );
buf ( n2326 , n204 );
buf ( n2327 , n2326 );
buf ( n2328 , n203 );
buf ( n2329 , n2328 );
buf ( n2330 , n202 );
buf ( n2331 , n2330 );
buf ( n2332 , n201 );
buf ( n2333 , n2332 );
buf ( n2334 , n200 );
buf ( n2335 , n2334 );
buf ( n2336 , n199 );
buf ( n2337 , n2336 );
buf ( n2338 , n198 );
buf ( n2339 , n2338 );
buf ( n2340 , n197 );
buf ( n2341 , n2340 );
buf ( n2342 , n196 );
buf ( n2343 , n2342 );
buf ( n2344 , n195 );
buf ( n2345 , n2344 );
buf ( n2346 , n194 );
buf ( n2347 , n2346 );
buf ( n2348 , n193 );
buf ( n2349 , n2348 );
buf ( n2350 , n192 );
buf ( n2351 , n2350 );
buf ( n2352 , n191 );
buf ( n2353 , n2352 );
buf ( n2354 , n242 );
buf ( n2355 , n2354 );
buf ( n2356 , n241 );
buf ( n2357 , n2356 );
buf ( n2358 , n240 );
buf ( n2359 , n2358 );
buf ( n2360 , n239 );
buf ( n2361 , n2360 );
buf ( n2362 , n238 );
buf ( n2363 , n2362 );
buf ( n2364 , n237 );
buf ( n2365 , n2364 );
buf ( n2366 , n236 );
buf ( n2367 , n2366 );
buf ( n2368 , n235 );
buf ( n2369 , n2368 );
buf ( n2370 , n234 );
buf ( n2371 , n2370 );
buf ( n2372 , n233 );
buf ( n2373 , n2372 );
buf ( n2374 , n232 );
buf ( n2375 , n2374 );
buf ( n2376 , n231 );
buf ( n2377 , n2376 );
buf ( n2378 , n230 );
buf ( n2379 , n2378 );
buf ( n2380 , n229 );
buf ( n2381 , n2380 );
buf ( n2382 , n228 );
buf ( n2383 , n2382 );
buf ( n2384 , n227 );
buf ( n2385 , n2384 );
buf ( n2386 , n226 );
buf ( n2387 , n2386 );
buf ( n2388 , n225 );
buf ( n2389 , n2388 );
buf ( n2390 , n224 );
buf ( n2391 , n2390 );
buf ( n2392 , n223 );
buf ( n2393 , n2392 );
buf ( n2394 , n222 );
buf ( n2395 , n2394 );
buf ( n2396 , n221 );
buf ( n2397 , n2396 );
buf ( n2398 , n220 );
buf ( n2399 , n2398 );
buf ( n2400 , n219 );
buf ( n2401 , n2400 );
buf ( n2402 , n218 );
buf ( n2403 , n2402 );
buf ( n2404 , n217 );
buf ( n2405 , n2404 );
buf ( n2406 , n216 );
buf ( n2407 , n2406 );
buf ( n2408 , n215 );
buf ( n2409 , n2408 );
buf ( n2410 , n214 );
buf ( n2411 , n2410 );
buf ( n2412 , n213 );
buf ( n2413 , n2412 );
buf ( n2414 , n212 );
buf ( n2415 , n2414 );
buf ( n2416 , n211 );
buf ( n2417 , n2416 );
buf ( n2418 , DFF_rd_reg_Q );
buf ( n2419 , n2418 );
buf ( n2420 , DFF_wr_reg_Q );
buf ( n2421 , n2420 );
buf ( n2422 , DFF_state_reg_Q );
not ( n2423 , n2282 );
and ( n2424 , n2282 , n2423 );
buf ( n2425 , n2424 );
buf ( n2426 , n2281 );
buf ( n2427 , n2280 );
not ( n2428 , n2422 );
buf ( n2429 , n2428 );
buf ( n2430 , n32 );
buf ( n2431 , n2424 );
buf ( n2432 , n2281 );
buf ( n2433 , n2280 );
and ( n2434 , n2430 , n2422 );
and ( n2435 , n2313 , n2428 );
or ( n2436 , n2434 , n2435 );
buf ( n2437 , n2436 );
buf ( n2438 , n33 );
buf ( n2439 , n2424 );
buf ( n2440 , n2281 );
buf ( n2441 , n2280 );
buf ( n2442 , n63 );
not ( n2443 , n2442 );
and ( n2444 , n2443 , n2438 );
not ( n2445 , n2438 );
not ( n2446 , n2430 );
xor ( n2447 , n2445 , n2446 );
and ( n2448 , n2447 , n2442 );
or ( n2449 , n2444 , n2448 );
and ( n2450 , n2449 , n2422 );
and ( n2451 , n2312 , n2428 );
or ( n2452 , n2450 , n2451 );
buf ( n2453 , n2452 );
buf ( n2454 , n34 );
buf ( n2455 , n2424 );
buf ( n2456 , n2281 );
buf ( n2457 , n2280 );
not ( n2458 , n2442 );
and ( n2459 , n2458 , n2454 );
not ( n2460 , n2454 );
and ( n2461 , n2445 , n2446 );
xor ( n2462 , n2460 , n2461 );
and ( n2463 , n2462 , n2442 );
or ( n2464 , n2459 , n2463 );
and ( n2465 , n2464 , n2422 );
and ( n2466 , n2311 , n2428 );
xor ( n2467 , n2465 , n2466 );
buf ( n2468 , n2467 );
buf ( n2469 , n35 );
buf ( n2470 , n2424 );
buf ( n2471 , n2281 );
buf ( n2472 , n2280 );
not ( n2473 , n2442 );
and ( n2474 , n2473 , n2469 );
not ( n2475 , n2469 );
and ( n2476 , n2460 , n2461 );
xor ( n2477 , n2475 , n2476 );
and ( n2478 , n2477 , n2442 );
or ( n2479 , n2474 , n2478 );
and ( n2480 , n2479 , n2422 );
and ( n2481 , n2310 , n2428 );
or ( n2482 , n2480 , n2481 );
buf ( n2483 , n2482 );
buf ( n2484 , n36 );
buf ( n2485 , n2424 );
buf ( n2486 , n2281 );
buf ( n2487 , n2280 );
not ( n2488 , n2442 );
and ( n2489 , n2488 , n2484 );
not ( n2490 , n2484 );
and ( n2491 , n2475 , n2476 );
xor ( n2492 , n2490 , n2491 );
and ( n2493 , n2492 , n2442 );
or ( n2494 , n2489 , n2493 );
and ( n2495 , n2494 , n2422 );
and ( n2496 , n2309 , n2428 );
or ( n2497 , n2495 , n2496 );
buf ( n2498 , n2497 );
buf ( n2499 , n37 );
buf ( n2500 , n2424 );
buf ( n2501 , n2281 );
buf ( n2502 , n2280 );
not ( n2503 , n2442 );
and ( n2504 , n2503 , n2499 );
not ( n2505 , n2499 );
and ( n2506 , n2490 , n2491 );
xor ( n2507 , n2505 , n2506 );
and ( n2508 , n2507 , n2442 );
or ( n2509 , n2504 , n2508 );
and ( n2510 , n2509 , n2422 );
and ( n2511 , n2308 , n2428 );
or ( n2512 , n2510 , n2511 );
buf ( n2513 , n2512 );
buf ( n2514 , n38 );
buf ( n2515 , n2424 );
buf ( n2516 , n2281 );
buf ( n2517 , n2280 );
not ( n2518 , n2442 );
and ( n2519 , n2518 , n2514 );
not ( n2520 , n2514 );
and ( n2521 , n2505 , n2506 );
xor ( n2522 , n2520 , n2521 );
and ( n2523 , n2522 , n2442 );
or ( n2524 , n2519 , n2523 );
and ( n2525 , n2524 , n2422 );
and ( n2526 , n2307 , n2428 );
or ( n2527 , n2525 , n2526 );
buf ( n2528 , n2527 );
buf ( n2529 , n39 );
buf ( n2530 , n2424 );
buf ( n2531 , n2281 );
buf ( n2532 , n2280 );
not ( n2533 , n2442 );
and ( n2534 , n2533 , n2529 );
not ( n2535 , n2529 );
and ( n2536 , n2520 , n2521 );
xor ( n2537 , n2535 , n2536 );
and ( n2538 , n2537 , n2442 );
or ( n2539 , n2534 , n2538 );
and ( n2540 , n2539 , n2422 );
and ( n2541 , n2306 , n2428 );
or ( n2542 , n2540 , n2541 );
buf ( n2543 , n2542 );
buf ( n2544 , n40 );
buf ( n2545 , n2424 );
buf ( n2546 , n2281 );
buf ( n2547 , n2280 );
not ( n2548 , n2442 );
and ( n2549 , n2548 , n2544 );
not ( n2550 , n2544 );
and ( n2551 , n2535 , n2536 );
xor ( n2552 , n2550 , n2551 );
and ( n2553 , n2552 , n2442 );
or ( n2554 , n2549 , n2553 );
and ( n2555 , n2554 , n2422 );
and ( n2556 , n2305 , n2428 );
or ( n2557 , n2555 , n2556 );
buf ( n2558 , n2557 );
buf ( n2559 , n41 );
buf ( n2560 , n2424 );
buf ( n2561 , n2281 );
buf ( n2562 , n2280 );
not ( n2563 , n2442 );
and ( n2564 , n2563 , n2559 );
not ( n2565 , n2559 );
and ( n2566 , n2550 , n2551 );
xor ( n2567 , n2565 , n2566 );
and ( n2568 , n2567 , n2442 );
or ( n2569 , n2564 , n2568 );
and ( n2570 , n2569 , n2422 );
and ( n2571 , n2304 , n2428 );
or ( n2572 , n2570 , n2571 );
buf ( n2573 , n2572 );
buf ( n2574 , n42 );
buf ( n2575 , n2424 );
buf ( n2576 , n2281 );
buf ( n2577 , n2280 );
not ( n2578 , n2442 );
and ( n2579 , n2578 , n2574 );
not ( n2580 , n2574 );
and ( n2581 , n2565 , n2566 );
xor ( n2582 , n2580 , n2581 );
and ( n2583 , n2582 , n2442 );
or ( n2584 , n2579 , n2583 );
and ( n2585 , n2584 , n2422 );
and ( n2586 , n2303 , n2428 );
or ( n2587 , n2585 , n2586 );
buf ( n2588 , n2587 );
buf ( n2589 , n43 );
buf ( n2590 , n2424 );
buf ( n2591 , n2281 );
buf ( n2592 , n2280 );
not ( n2593 , n2442 );
and ( n2594 , n2593 , n2589 );
not ( n2595 , n2589 );
and ( n2596 , n2580 , n2581 );
xor ( n2597 , n2595 , n2596 );
and ( n2598 , n2597 , n2442 );
or ( n2599 , n2594 , n2598 );
and ( n2600 , n2599 , n2422 );
and ( n2601 , n2302 , n2428 );
or ( n2602 , n2600 , n2601 );
buf ( n2603 , n2602 );
buf ( n2604 , n44 );
buf ( n2605 , n2424 );
buf ( n2606 , n2281 );
buf ( n2607 , n2280 );
not ( n2608 , n2442 );
and ( n2609 , n2608 , n2604 );
not ( n2610 , n2604 );
and ( n2611 , n2595 , n2596 );
xor ( n2612 , n2610 , n2611 );
and ( n2613 , n2612 , n2442 );
or ( n2614 , n2609 , n2613 );
and ( n2615 , n2614 , n2422 );
and ( n2616 , n2301 , n2428 );
or ( n2617 , n2615 , n2616 );
buf ( n2618 , n2617 );
buf ( n2619 , n45 );
buf ( n2620 , n2424 );
buf ( n2621 , n2281 );
buf ( n2622 , n2280 );
not ( n2623 , n2442 );
and ( n2624 , n2623 , n2619 );
not ( n2625 , n2619 );
and ( n2626 , n2610 , n2611 );
xor ( n2627 , n2625 , n2626 );
and ( n2628 , n2627 , n2442 );
or ( n2629 , n2624 , n2628 );
and ( n2630 , n2629 , n2422 );
and ( n2631 , n2300 , n2428 );
or ( n2632 , n2630 , n2631 );
buf ( n2633 , n2632 );
buf ( n2634 , n46 );
buf ( n2635 , n2424 );
buf ( n2636 , n2281 );
buf ( n2637 , n2280 );
not ( n2638 , n2442 );
and ( n2639 , n2638 , n2634 );
not ( n2640 , n2634 );
and ( n2641 , n2625 , n2626 );
xor ( n2642 , n2640 , n2641 );
and ( n2643 , n2642 , n2442 );
or ( n2644 , n2639 , n2643 );
and ( n2645 , n2644 , n2422 );
and ( n2646 , n2299 , n2428 );
or ( n2647 , n2645 , n2646 );
buf ( n2648 , n2647 );
buf ( n2649 , n47 );
buf ( n2650 , n2424 );
buf ( n2651 , n2281 );
buf ( n2652 , n2280 );
not ( n2653 , n2442 );
and ( n2654 , n2653 , n2649 );
not ( n2655 , n2649 );
and ( n2656 , n2640 , n2641 );
xor ( n2657 , n2655 , n2656 );
and ( n2658 , n2657 , n2442 );
or ( n2659 , n2654 , n2658 );
and ( n2660 , n2659 , n2422 );
and ( n2661 , n2298 , n2428 );
or ( n2662 , n2660 , n2661 );
buf ( n2663 , n2662 );
buf ( n2664 , n48 );
buf ( n2665 , n2424 );
buf ( n2666 , n2281 );
buf ( n2667 , n2280 );
not ( n2668 , n2442 );
and ( n2669 , n2668 , n2664 );
not ( n2670 , n2664 );
and ( n2671 , n2655 , n2656 );
xor ( n2672 , n2670 , n2671 );
and ( n2673 , n2672 , n2442 );
or ( n2674 , n2669 , n2673 );
and ( n2675 , n2674 , n2422 );
and ( n2676 , n2297 , n2428 );
or ( n2677 , n2675 , n2676 );
buf ( n2678 , n2677 );
buf ( n2679 , n49 );
buf ( n2680 , n2424 );
buf ( n2681 , n2281 );
buf ( n2682 , n2280 );
not ( n2683 , n2442 );
and ( n2684 , n2683 , n2679 );
not ( n2685 , n2679 );
and ( n2686 , n2670 , n2671 );
xor ( n2687 , n2685 , n2686 );
and ( n2688 , n2687 , n2442 );
or ( n2689 , n2684 , n2688 );
and ( n2690 , n2689 , n2422 );
and ( n2691 , n2296 , n2428 );
or ( n2692 , n2690 , n2691 );
buf ( n2693 , n2692 );
buf ( n2694 , n50 );
buf ( n2695 , n2424 );
buf ( n2696 , n2281 );
buf ( n2697 , n2280 );
not ( n2698 , n2442 );
and ( n2699 , n2698 , n2694 );
not ( n2700 , n2694 );
and ( n2701 , n2685 , n2686 );
xor ( n2702 , n2700 , n2701 );
and ( n2703 , n2702 , n2442 );
or ( n2704 , n2699 , n2703 );
and ( n2705 , n2704 , n2422 );
and ( n2706 , n2295 , n2428 );
or ( n2707 , n2705 , n2706 );
buf ( n2708 , n2707 );
buf ( n2709 , n51 );
buf ( n2710 , n2424 );
buf ( n2711 , n2281 );
buf ( n2712 , n2280 );
not ( n2713 , n2442 );
and ( n2714 , n2713 , n2709 );
not ( n2715 , n2709 );
and ( n2716 , n2700 , n2701 );
xor ( n2717 , n2715 , n2716 );
and ( n2718 , n2717 , n2442 );
or ( n2719 , n2714 , n2718 );
and ( n2720 , n2719 , n2422 );
and ( n2721 , n2294 , n2428 );
or ( n2722 , n2720 , n2721 );
buf ( n2723 , n2722 );
buf ( n2724 , n52 );
buf ( n2725 , n2424 );
buf ( n2726 , n2281 );
buf ( n2727 , n2280 );
not ( n2728 , n2442 );
and ( n2729 , n2728 , n2724 );
not ( n2730 , n2724 );
and ( n2731 , n2715 , n2716 );
xor ( n2732 , n2730 , n2731 );
and ( n2733 , n2732 , n2442 );
or ( n2734 , n2729 , n2733 );
and ( n2735 , n2734 , n2422 );
and ( n2736 , n2293 , n2428 );
or ( n2737 , n2735 , n2736 );
buf ( n2738 , n2737 );
buf ( n2739 , n53 );
buf ( n2740 , n2424 );
buf ( n2741 , n2281 );
buf ( n2742 , n2280 );
not ( n2743 , n2442 );
and ( n2744 , n2743 , n2739 );
not ( n2745 , n2739 );
and ( n2746 , n2730 , n2731 );
xor ( n2747 , n2745 , n2746 );
and ( n2748 , n2747 , n2442 );
or ( n2749 , n2744 , n2748 );
and ( n2750 , n2749 , n2422 );
and ( n2751 , n2292 , n2428 );
or ( n2752 , n2750 , n2751 );
buf ( n2753 , n2752 );
buf ( n2754 , n54 );
buf ( n2755 , n2424 );
buf ( n2756 , n2281 );
buf ( n2757 , n2280 );
not ( n2758 , n2442 );
and ( n2759 , n2758 , n2754 );
not ( n2760 , n2754 );
and ( n2761 , n2745 , n2746 );
xor ( n2762 , n2760 , n2761 );
and ( n2763 , n2762 , n2442 );
or ( n2764 , n2759 , n2763 );
and ( n2765 , n2764 , n2422 );
and ( n2766 , n2291 , n2428 );
or ( n2767 , n2765 , n2766 );
buf ( n2768 , n2767 );
buf ( n2769 , n55 );
buf ( n2770 , n2424 );
buf ( n2771 , n2281 );
buf ( n2772 , n2280 );
not ( n2773 , n2442 );
and ( n2774 , n2773 , n2769 );
not ( n2775 , n2769 );
and ( n2776 , n2760 , n2761 );
xor ( n2777 , n2775 , n2776 );
and ( n2778 , n2777 , n2442 );
or ( n2779 , n2774 , n2778 );
and ( n2780 , n2779 , n2422 );
and ( n2781 , n2290 , n2428 );
or ( n2782 , n2780 , n2781 );
buf ( n2783 , n2782 );
buf ( n2784 , n56 );
buf ( n2785 , n2424 );
buf ( n2786 , n2281 );
buf ( n2787 , n2280 );
not ( n2788 , n2442 );
and ( n2789 , n2788 , n2784 );
not ( n2790 , n2784 );
and ( n2791 , n2775 , n2776 );
xor ( n2792 , n2790 , n2791 );
and ( n2793 , n2792 , n2442 );
or ( n2794 , n2789 , n2793 );
and ( n2795 , n2794 , n2422 );
and ( n2796 , n2289 , n2428 );
or ( n2797 , n2795 , n2796 );
buf ( n2798 , n2797 );
buf ( n2799 , n57 );
buf ( n2800 , n2424 );
buf ( n2801 , n2281 );
buf ( n2802 , n2280 );
not ( n2803 , n2442 );
and ( n2804 , n2803 , n2799 );
not ( n2805 , n2799 );
and ( n2806 , n2790 , n2791 );
xor ( n2807 , n2805 , n2806 );
and ( n2808 , n2807 , n2442 );
or ( n2809 , n2804 , n2808 );
and ( n2810 , n2809 , n2422 );
and ( n2811 , n2288 , n2428 );
or ( n2812 , n2810 , n2811 );
buf ( n2813 , n2812 );
buf ( n2814 , n58 );
buf ( n2815 , n2424 );
buf ( n2816 , n2281 );
buf ( n2817 , n2280 );
not ( n2818 , n2442 );
and ( n2819 , n2818 , n2814 );
not ( n2820 , n2814 );
and ( n2821 , n2805 , n2806 );
xor ( n2822 , n2820 , n2821 );
and ( n2823 , n2822 , n2442 );
or ( n2824 , n2819 , n2823 );
and ( n2825 , n2824 , n2422 );
and ( n2826 , n2287 , n2428 );
or ( n2827 , n2825 , n2826 );
buf ( n2828 , n2827 );
buf ( n2829 , n59 );
buf ( n2830 , n2424 );
buf ( n2831 , n2281 );
buf ( n2832 , n2280 );
not ( n2833 , n2442 );
and ( n2834 , n2833 , n2829 );
not ( n2835 , n2829 );
and ( n2836 , n2820 , n2821 );
xor ( n2837 , n2835 , n2836 );
and ( n2838 , n2837 , n2442 );
or ( n2839 , n2834 , n2838 );
and ( n2840 , n2839 , n2422 );
and ( n2841 , n2286 , n2428 );
or ( n2842 , n2840 , n2841 );
buf ( n2843 , n2842 );
buf ( n2844 , n60 );
buf ( n2845 , n2424 );
buf ( n2846 , n2281 );
buf ( n2847 , n2280 );
not ( n2848 , n2442 );
and ( n2849 , n2848 , n2844 );
not ( n2850 , n2844 );
and ( n2851 , n2835 , n2836 );
xor ( n2852 , n2850 , n2851 );
and ( n2853 , n2852 , n2442 );
or ( n2854 , n2849 , n2853 );
and ( n2855 , n2854 , n2422 );
and ( n2856 , n2285 , n2428 );
or ( n2857 , n2855 , n2856 );
buf ( n2858 , n2857 );
buf ( n2859 , n61 );
buf ( n2860 , n2424 );
buf ( n2861 , n2281 );
buf ( n2862 , n2280 );
not ( n2863 , n2442 );
and ( n2864 , n2863 , n2859 );
not ( n2865 , n2859 );
and ( n2866 , n2850 , n2851 );
xor ( n2867 , n2865 , n2866 );
and ( n2868 , n2867 , n2442 );
or ( n2869 , n2864 , n2868 );
and ( n2870 , n2869 , n2422 );
and ( n2871 , n2284 , n2428 );
or ( n2872 , n2870 , n2871 );
buf ( n2873 , n2872 );
buf ( n2874 , n62 );
buf ( n2875 , n2424 );
buf ( n2876 , n2281 );
buf ( n2877 , n2280 );
not ( n2878 , n2442 );
and ( n2879 , n2878 , n2874 );
not ( n2880 , n2874 );
and ( n2881 , n2865 , n2866 );
xor ( n2882 , n2880 , n2881 );
and ( n2883 , n2882 , n2442 );
or ( n2884 , n2879 , n2883 );
and ( n2885 , n2884 , n2422 );
and ( n2886 , n2283 , n2428 );
or ( n2887 , n2885 , n2886 );
buf ( n2888 , n2887 );
buf ( n2889 , n2424 );
buf ( n2890 , n2281 );
buf ( n2891 , n2280 );
buf ( n2892 , n2442 );
not ( n2893 , n2892 );
and ( n2894 , n2893 , n2442 );
not ( n2895 , n2442 );
and ( n2896 , n2880 , n2881 );
xor ( n2897 , n2895 , n2896 );
and ( n2898 , n2897 , n2892 );
or ( n2899 , n2894 , n2898 );
and ( n2900 , n2899 , n2422 );
and ( n2901 , n2282 , n2428 );
or ( n2902 , n2900 , n2901 );
buf ( n2903 , n2902 );
buf ( n2904 , n64 );
buf ( n2905 , n2424 );
buf ( n2906 , n2281 );
buf ( n2907 , n2280 );
not ( n2908 , n2899 );
and ( n2909 , n2908 , n2779 );
not ( n2910 , n2779 );
not ( n2911 , n2764 );
not ( n2912 , n2749 );
not ( n2913 , n2734 );
not ( n2914 , n2719 );
not ( n2915 , n2704 );
not ( n2916 , n2689 );
not ( n2917 , n2674 );
not ( n2918 , n2659 );
not ( n2919 , n2644 );
not ( n2920 , n2629 );
not ( n2921 , n2614 );
not ( n2922 , n2599 );
not ( n2923 , n2584 );
not ( n2924 , n2569 );
not ( n2925 , n2554 );
not ( n2926 , n2539 );
not ( n2927 , n2524 );
not ( n2928 , n2509 );
not ( n2929 , n2494 );
not ( n2930 , n2479 );
not ( n2931 , n2464 );
not ( n2932 , n2449 );
not ( n2933 , n2430 );
nand ( n2934 , n2932 , n2933 );
and ( n2935 , n2931 , n2934 );
and ( n2936 , n2930 , n2935 );
and ( n2937 , n2929 , n2936 );
and ( n2938 , n2928 , n2937 );
and ( n2939 , n2927 , n2938 );
and ( n2940 , n2926 , n2939 );
and ( n2941 , n2925 , n2940 );
and ( n2942 , n2924 , n2941 );
and ( n2943 , n2923 , n2942 );
and ( n2944 , n2922 , n2943 );
and ( n2945 , n2921 , n2944 );
and ( n2946 , n2920 , n2945 );
and ( n2947 , n2919 , n2946 );
and ( n2948 , n2918 , n2947 );
and ( n2949 , n2917 , n2948 );
and ( n2950 , n2916 , n2949 );
and ( n2951 , n2915 , n2950 );
and ( n2952 , n2914 , n2951 );
and ( n2953 , n2913 , n2952 );
and ( n2954 , n2912 , n2953 );
and ( n2955 , n2911 , n2954 );
xor ( n2956 , n2910 , n2955 );
and ( n2957 , n2956 , n2899 );
or ( n2958 , n2909 , n2957 );
not ( n2959 , n2958 );
not ( n2960 , n2959 );
not ( n2961 , n2960 );
not ( n2962 , n2961 );
buf ( n2963 , n2962 );
buf ( n2964 , n2963 );
not ( n2965 , n2899 );
and ( n2966 , n2965 , n2424 );
buf ( n2967 , n2899 );
not ( n2968 , n2967 );
and ( n2969 , n2968 , n2899 );
not ( n2970 , n2899 );
not ( n2971 , n2884 );
not ( n2972 , n2869 );
not ( n2973 , n2854 );
not ( n2974 , n2839 );
not ( n2975 , n2824 );
not ( n2976 , n2809 );
not ( n2977 , n2794 );
and ( n2978 , n2910 , n2955 );
and ( n2979 , n2977 , n2978 );
and ( n2980 , n2976 , n2979 );
and ( n2981 , n2975 , n2980 );
and ( n2982 , n2974 , n2981 );
and ( n2983 , n2973 , n2982 );
and ( n2984 , n2972 , n2983 );
and ( n2985 , n2971 , n2984 );
xor ( n2986 , n2970 , n2985 );
and ( n2987 , n2986 , n2967 );
or ( n2988 , n2969 , n2987 );
not ( n2989 , n2988 );
not ( n2990 , n2989 );
not ( n2991 , n2990 );
not ( n2992 , n2899 );
and ( n2993 , n2992 , n2884 );
xor ( n2994 , n2971 , n2984 );
and ( n2995 , n2994 , n2899 );
or ( n2996 , n2993 , n2995 );
not ( n2997 , n2996 );
not ( n2998 , n2997 );
not ( n2999 , n2998 );
not ( n3000 , n2899 );
and ( n3001 , n3000 , n2869 );
xor ( n3002 , n2972 , n2983 );
and ( n3003 , n3002 , n2899 );
or ( n3004 , n3001 , n3003 );
not ( n3005 , n3004 );
not ( n3006 , n3005 );
not ( n3007 , n3006 );
not ( n3008 , n2899 );
and ( n3009 , n3008 , n2854 );
xor ( n3010 , n2973 , n2982 );
and ( n3011 , n3010 , n2899 );
or ( n3012 , n3009 , n3011 );
not ( n3013 , n3012 );
not ( n3014 , n3013 );
not ( n3015 , n3014 );
not ( n3016 , n2899 );
and ( n3017 , n3016 , n2839 );
xor ( n3018 , n2974 , n2981 );
and ( n3019 , n3018 , n2899 );
or ( n3020 , n3017 , n3019 );
not ( n3021 , n3020 );
not ( n3022 , n3021 );
not ( n3023 , n3022 );
not ( n3024 , n2899 );
and ( n3025 , n3024 , n2824 );
xor ( n3026 , n2975 , n2980 );
and ( n3027 , n3026 , n2899 );
or ( n3028 , n3025 , n3027 );
not ( n3029 , n3028 );
not ( n3030 , n3029 );
not ( n3031 , n3030 );
not ( n3032 , n2899 );
and ( n3033 , n3032 , n2809 );
xor ( n3034 , n2976 , n2979 );
and ( n3035 , n3034 , n2899 );
or ( n3036 , n3033 , n3035 );
not ( n3037 , n3036 );
not ( n3038 , n3037 );
not ( n3039 , n3038 );
not ( n3040 , n2899 );
and ( n3041 , n3040 , n2794 );
xor ( n3042 , n2977 , n2978 );
and ( n3043 , n3042 , n2899 );
or ( n3044 , n3041 , n3043 );
not ( n3045 , n3044 );
not ( n3046 , n3045 );
not ( n3047 , n3046 );
not ( n3048 , n2960 );
and ( n3049 , n3047 , n3048 );
and ( n3050 , n3039 , n3049 );
and ( n3051 , n3031 , n3050 );
and ( n3052 , n3023 , n3051 );
and ( n3053 , n3015 , n3052 );
and ( n3054 , n3007 , n3053 );
and ( n3055 , n2999 , n3054 );
and ( n3056 , n2991 , n3055 );
not ( n3057 , n3056 );
and ( n3058 , n3057 , n2899 );
or ( n3059 , n2966 , n3058 );
and ( n3060 , n2964 , n3059 );
not ( n3061 , n3060 );
and ( n3062 , n3061 , n2962 );
xor ( n3063 , n2962 , n3059 );
xor ( n3064 , n3063 , n3059 );
and ( n3065 , n3064 , n3060 );
or ( n3066 , n3062 , n3065 );
not ( n3067 , n2899 );
and ( n3068 , n3067 , n2794 );
not ( n3069 , n2794 );
not ( n3070 , n2779 );
not ( n3071 , n2764 );
not ( n3072 , n2749 );
not ( n3073 , n2734 );
not ( n3074 , n2719 );
not ( n3075 , n2704 );
not ( n3076 , n2689 );
not ( n3077 , n2674 );
not ( n3078 , n2659 );
not ( n3079 , n2644 );
not ( n3080 , n2629 );
not ( n3081 , n2614 );
not ( n3082 , n2599 );
not ( n3083 , n2584 );
not ( n3084 , n2569 );
not ( n3085 , n2554 );
not ( n3086 , n2539 );
not ( n3087 , n2524 );
not ( n3088 , n2509 );
not ( n3089 , n2494 );
not ( n3090 , n2479 );
not ( n3091 , n2464 );
not ( n3092 , n2449 );
not ( n3093 , n2430 );
and ( n3094 , n3092 , n3093 );
and ( n3095 , n3091 , n3094 );
and ( n3096 , n3090 , n3095 );
and ( n3097 , n3089 , n3096 );
and ( n3098 , n3088 , n3097 );
and ( n3099 , n3087 , n3098 );
and ( n3100 , n3086 , n3099 );
and ( n3101 , n3085 , n3100 );
and ( n3102 , n3084 , n3101 );
and ( n3103 , n3083 , n3102 );
and ( n3104 , n3082 , n3103 );
and ( n3105 , n3081 , n3104 );
and ( n3106 , n3080 , n3105 );
and ( n3107 , n3079 , n3106 );
and ( n3108 , n3078 , n3107 );
and ( n3109 , n3077 , n3108 );
and ( n3110 , n3076 , n3109 );
and ( n3111 , n3075 , n3110 );
and ( n3112 , n3074 , n3111 );
and ( n3113 , n3073 , n3112 );
and ( n3114 , n3072 , n3113 );
and ( n3115 , n3071 , n3114 );
and ( n3116 , n3070 , n3115 );
xor ( n3117 , n3069 , n3116 );
and ( n3118 , n3117 , n2899 );
or ( n3119 , n3068 , n3118 );
not ( n3120 , n3119 );
not ( n3121 , n3120 );
not ( n3122 , n3121 );
not ( n3123 , n3122 );
not ( n3124 , n2899 );
and ( n3125 , n3124 , n2424 );
buf ( n3126 , n2899 );
not ( n3127 , n3126 );
and ( n3128 , n3127 , n2899 );
not ( n3129 , n2899 );
not ( n3130 , n2884 );
not ( n3131 , n2869 );
not ( n3132 , n2854 );
not ( n3133 , n2839 );
not ( n3134 , n2824 );
not ( n3135 , n2809 );
and ( n3136 , n3069 , n3116 );
and ( n3137 , n3135 , n3136 );
and ( n3138 , n3134 , n3137 );
and ( n3139 , n3133 , n3138 );
and ( n3140 , n3132 , n3139 );
and ( n3141 , n3131 , n3140 );
and ( n3142 , n3130 , n3141 );
xor ( n3143 , n3129 , n3142 );
and ( n3144 , n3143 , n3126 );
or ( n3145 , n3128 , n3144 );
not ( n3146 , n3145 );
not ( n3147 , n3146 );
not ( n3148 , n3147 );
not ( n3149 , n2899 );
and ( n3150 , n3149 , n2884 );
xor ( n3151 , n3130 , n3141 );
and ( n3152 , n3151 , n2899 );
or ( n3153 , n3150 , n3152 );
not ( n3154 , n3153 );
not ( n3155 , n3154 );
not ( n3156 , n3155 );
not ( n3157 , n2899 );
and ( n3158 , n3157 , n2869 );
xor ( n3159 , n3131 , n3140 );
and ( n3160 , n3159 , n2899 );
or ( n3161 , n3158 , n3160 );
not ( n3162 , n3161 );
not ( n3163 , n3162 );
not ( n3164 , n3163 );
not ( n3165 , n2899 );
and ( n3166 , n3165 , n2854 );
xor ( n3167 , n3132 , n3139 );
and ( n3168 , n3167 , n2899 );
or ( n3169 , n3166 , n3168 );
not ( n3170 , n3169 );
not ( n3171 , n3170 );
not ( n3172 , n3171 );
not ( n3173 , n2899 );
and ( n3174 , n3173 , n2839 );
xor ( n3175 , n3133 , n3138 );
and ( n3176 , n3175 , n2899 );
or ( n3177 , n3174 , n3176 );
not ( n3178 , n3177 );
not ( n3179 , n3178 );
not ( n3180 , n3179 );
not ( n3181 , n2899 );
and ( n3182 , n3181 , n2824 );
xor ( n3183 , n3134 , n3137 );
and ( n3184 , n3183 , n2899 );
or ( n3185 , n3182 , n3184 );
not ( n3186 , n3185 );
not ( n3187 , n3186 );
not ( n3188 , n3187 );
not ( n3189 , n2899 );
and ( n3190 , n3189 , n2809 );
xor ( n3191 , n3135 , n3136 );
and ( n3192 , n3191 , n2899 );
or ( n3193 , n3190 , n3192 );
not ( n3194 , n3193 );
not ( n3195 , n3194 );
not ( n3196 , n3195 );
not ( n3197 , n3121 );
and ( n3198 , n3196 , n3197 );
and ( n3199 , n3188 , n3198 );
and ( n3200 , n3180 , n3199 );
and ( n3201 , n3172 , n3200 );
and ( n3202 , n3164 , n3201 );
and ( n3203 , n3156 , n3202 );
and ( n3204 , n3148 , n3203 );
not ( n3205 , n3204 );
and ( n3206 , n3205 , n2899 );
or ( n3207 , n3125 , n3206 );
not ( n3208 , n3207 );
not ( n3209 , n2899 );
and ( n3210 , n3209 , n3195 );
xor ( n3211 , n3196 , n3197 );
and ( n3212 , n3211 , n2899 );
or ( n3213 , n3210 , n3212 );
and ( n3214 , n3208 , n3213 );
not ( n3215 , n3213 );
not ( n3216 , n3121 );
xor ( n3217 , n3215 , n3216 );
and ( n3218 , n3217 , n3207 );
or ( n3219 , n3214 , n3218 );
not ( n3220 , n3219 );
not ( n3221 , n3220 );
or ( n3222 , n3123 , n3221 );
not ( n3223 , n3207 );
not ( n3224 , n2899 );
and ( n3225 , n3224 , n3187 );
xor ( n3226 , n3188 , n3198 );
and ( n3227 , n3226 , n2899 );
or ( n3228 , n3225 , n3227 );
and ( n3229 , n3223 , n3228 );
not ( n3230 , n3228 );
and ( n3231 , n3215 , n3216 );
xor ( n3232 , n3230 , n3231 );
and ( n3233 , n3232 , n3207 );
or ( n3234 , n3229 , n3233 );
not ( n3235 , n3234 );
not ( n3236 , n3235 );
or ( n3237 , n3222 , n3236 );
and ( n3238 , n3237 , n3207 );
not ( n3239 , n3238 );
and ( n3240 , n3239 , n3123 );
xor ( n3241 , n3123 , n3207 );
xor ( n3242 , n3241 , n3207 );
and ( n3243 , n3242 , n3238 );
or ( n3244 , n3240 , n3243 );
not ( n3245 , n3238 );
and ( n3246 , n3245 , n3221 );
xor ( n3247 , n3221 , n3207 );
and ( n3248 , n3241 , n3207 );
xor ( n3249 , n3247 , n3248 );
and ( n3250 , n3249 , n3238 );
or ( n3251 , n3246 , n3250 );
not ( n3252 , n3238 );
and ( n3253 , n3252 , n3236 );
xor ( n3254 , n3236 , n3207 );
and ( n3255 , n3247 , n3248 );
xor ( n3256 , n3254 , n3255 );
and ( n3257 , n3256 , n3238 );
or ( n3258 , n3253 , n3257 );
and ( n3259 , n3244 , n3251 , n3258 );
or ( n3260 , n3066 , n3259 );
not ( n3261 , n3260 );
not ( n3262 , n3244 );
not ( n3263 , n3258 );
nor ( n3264 , n3262 , n3251 , n3263 );
not ( n3265 , n3264 );
nor ( n3266 , n3244 , n3251 , n3263 );
not ( n3267 , n3266 );
and ( n3268 , n3244 , n3251 , n3263 );
not ( n3269 , n3268 );
and ( n3270 , n3262 , n3251 , n3263 );
not ( n3271 , n3270 );
nor ( n3272 , n3262 , n3251 , n3258 );
not ( n3273 , n3272 );
nor ( n3274 , n3244 , n3251 , n3258 );
not ( n3275 , n3274 );
and ( n3276 , n3275 , n2904 );
and ( n3277 , n2424 , n3274 );
or ( n3278 , n3276 , n3277 );
and ( n3279 , n3273 , n3278 );
or ( n3280 , n2282 , n2423 );
and ( n3281 , n3280 , n3272 );
or ( n3282 , n3279 , n3281 );
and ( n3283 , n3271 , n3282 );
and ( n3284 , n2424 , n3270 );
or ( n3285 , n3283 , n3284 );
and ( n3286 , n3269 , n3285 );
and ( n3287 , n3280 , n3268 );
or ( n3288 , n3286 , n3287 );
and ( n3289 , n3267 , n3288 );
buf ( n3290 , DFF_B_reg_Q );
not ( n3291 , n3290 );
and ( n3292 , n3291 , n2904 );
and ( n3293 , n3280 , n3290 );
or ( n3294 , n3292 , n3293 );
and ( n3295 , n3294 , n3266 );
or ( n3296 , n3289 , n3295 );
and ( n3297 , n3265 , n3296 );
not ( n3298 , n3290 );
not ( n3299 , n3298 );
and ( n3300 , n3299 , n2904 );
and ( n3301 , n3280 , n3298 );
or ( n3302 , n3300 , n3301 );
and ( n3303 , n3302 , n3264 );
or ( n3304 , n3297 , n3303 );
and ( n3305 , n3261 , n3304 );
and ( n3306 , n2904 , n3260 );
or ( n3307 , n3305 , n3306 );
and ( n3308 , n3307 , n2422 );
and ( n3309 , n2904 , n2428 );
or ( n3310 , n3308 , n3309 );
buf ( n3311 , n3310 );
buf ( n3312 , n65 );
buf ( n3313 , n2424 );
buf ( n3314 , n2281 );
buf ( n3315 , n2280 );
not ( n3316 , n3260 );
not ( n3317 , n3264 );
not ( n3318 , n3266 );
not ( n3319 , n3268 );
not ( n3320 , n3270 );
not ( n3321 , n3272 );
not ( n3322 , n3274 );
and ( n3323 , n3322 , n3312 );
and ( n3324 , n2424 , n3274 );
or ( n3325 , n3323 , n3324 );
and ( n3326 , n3321 , n3325 );
and ( n3327 , n2424 , n3272 );
or ( n3328 , n3326 , n3327 );
and ( n3329 , n3320 , n3328 );
and ( n3330 , n3280 , n3270 );
or ( n3331 , n3329 , n3330 );
and ( n3332 , n3319 , n3331 );
and ( n3333 , n3280 , n3268 );
or ( n3334 , n3332 , n3333 );
and ( n3335 , n3318 , n3334 );
not ( n3336 , n3290 );
and ( n3337 , n3336 , n3312 );
and ( n3338 , n3280 , n3290 );
or ( n3339 , n3337 , n3338 );
and ( n3340 , n3339 , n3266 );
or ( n3341 , n3335 , n3340 );
and ( n3342 , n3317 , n3341 );
not ( n3343 , n3298 );
and ( n3344 , n3343 , n3312 );
and ( n3345 , n3280 , n3298 );
or ( n3346 , n3344 , n3345 );
and ( n3347 , n3346 , n3264 );
or ( n3348 , n3342 , n3347 );
and ( n3349 , n3316 , n3348 );
and ( n3350 , n3312 , n3260 );
or ( n3351 , n3349 , n3350 );
and ( n3352 , n3351 , n2422 );
and ( n3353 , n3312 , n2428 );
or ( n3354 , n3352 , n3353 );
buf ( n3355 , n3354 );
buf ( n3356 , n66 );
buf ( n3357 , n2424 );
buf ( n3358 , n2281 );
buf ( n3359 , n2280 );
not ( n3360 , n3260 );
not ( n3361 , n3356 );
not ( n3362 , n3361 );
buf ( n3363 , n3362 );
not ( n3364 , n2899 );
and ( n3365 , n3364 , n2719 );
not ( n3366 , n2719 );
not ( n3367 , n2704 );
not ( n3368 , n2689 );
not ( n3369 , n2674 );
not ( n3370 , n2659 );
not ( n3371 , n2644 );
not ( n3372 , n2629 );
not ( n3373 , n2614 );
not ( n3374 , n2599 );
not ( n3375 , n2584 );
not ( n3376 , n2569 );
not ( n3377 , n2554 );
not ( n3378 , n2539 );
not ( n3379 , n2524 );
not ( n3380 , n2509 );
not ( n3381 , n2494 );
not ( n3382 , n2479 );
not ( n3383 , n2464 );
not ( n3384 , n2449 );
not ( n3385 , n2430 );
and ( n3386 , n3384 , n3385 );
and ( n3387 , n3383 , n3386 );
and ( n3388 , n3382 , n3387 );
and ( n3389 , n3381 , n3388 );
and ( n3390 , n3380 , n3389 );
and ( n3391 , n3379 , n3390 );
and ( n3392 , n3378 , n3391 );
and ( n3393 , n3377 , n3392 );
and ( n3394 , n3376 , n3393 );
and ( n3395 , n3375 , n3394 );
and ( n3396 , n3374 , n3395 );
and ( n3397 , n3373 , n3396 );
and ( n3398 , n3372 , n3397 );
and ( n3399 , n3371 , n3398 );
and ( n3400 , n3370 , n3399 );
and ( n3401 , n3369 , n3400 );
and ( n3402 , n3368 , n3401 );
and ( n3403 , n3367 , n3402 );
xor ( n3404 , n3366 , n3403 );
and ( n3405 , n3404 , n2899 );
or ( n3406 , n3365 , n3405 );
not ( n3407 , n3406 );
not ( n3408 , n3407 );
not ( n3409 , n3408 );
not ( n3410 , n3409 );
not ( n3411 , n2899 );
and ( n3412 , n3411 , n2424 );
buf ( n3413 , n2899 );
not ( n3414 , n3413 );
and ( n3415 , n3414 , n2899 );
not ( n3416 , n2899 );
not ( n3417 , n2884 );
not ( n3418 , n2869 );
not ( n3419 , n2854 );
not ( n3420 , n2839 );
not ( n3421 , n2824 );
not ( n3422 , n2809 );
not ( n3423 , n2794 );
not ( n3424 , n2779 );
not ( n3425 , n2764 );
not ( n3426 , n2749 );
not ( n3427 , n2734 );
and ( n3428 , n3366 , n3403 );
and ( n3429 , n3427 , n3428 );
and ( n3430 , n3426 , n3429 );
and ( n3431 , n3425 , n3430 );
and ( n3432 , n3424 , n3431 );
and ( n3433 , n3423 , n3432 );
and ( n3434 , n3422 , n3433 );
and ( n3435 , n3421 , n3434 );
and ( n3436 , n3420 , n3435 );
and ( n3437 , n3419 , n3436 );
and ( n3438 , n3418 , n3437 );
and ( n3439 , n3417 , n3438 );
xor ( n3440 , n3416 , n3439 );
and ( n3441 , n3440 , n3413 );
or ( n3442 , n3415 , n3441 );
not ( n3443 , n3442 );
not ( n3444 , n3443 );
not ( n3445 , n3444 );
not ( n3446 , n2899 );
and ( n3447 , n3446 , n2884 );
xor ( n3448 , n3417 , n3438 );
and ( n3449 , n3448 , n2899 );
or ( n3450 , n3447 , n3449 );
not ( n3451 , n3450 );
not ( n3452 , n3451 );
not ( n3453 , n3452 );
not ( n3454 , n2899 );
and ( n3455 , n3454 , n2869 );
xor ( n3456 , n3418 , n3437 );
and ( n3457 , n3456 , n2899 );
or ( n3458 , n3455 , n3457 );
not ( n3459 , n3458 );
not ( n3460 , n3459 );
not ( n3461 , n3460 );
not ( n3462 , n2899 );
and ( n3463 , n3462 , n2854 );
xor ( n3464 , n3419 , n3436 );
and ( n3465 , n3464 , n2899 );
or ( n3466 , n3463 , n3465 );
not ( n3467 , n3466 );
not ( n3468 , n3467 );
not ( n3469 , n3468 );
not ( n3470 , n2899 );
and ( n3471 , n3470 , n2839 );
xor ( n3472 , n3420 , n3435 );
and ( n3473 , n3472 , n2899 );
or ( n3474 , n3471 , n3473 );
not ( n3475 , n3474 );
not ( n3476 , n3475 );
not ( n3477 , n3476 );
not ( n3478 , n2899 );
and ( n3479 , n3478 , n2824 );
xor ( n3480 , n3421 , n3434 );
and ( n3481 , n3480 , n2899 );
or ( n3482 , n3479 , n3481 );
not ( n3483 , n3482 );
not ( n3484 , n3483 );
not ( n3485 , n3484 );
not ( n3486 , n2899 );
and ( n3487 , n3486 , n2809 );
xor ( n3488 , n3422 , n3433 );
and ( n3489 , n3488 , n2899 );
or ( n3490 , n3487 , n3489 );
not ( n3491 , n3490 );
not ( n3492 , n3491 );
not ( n3493 , n3492 );
not ( n3494 , n2899 );
and ( n3495 , n3494 , n2794 );
xor ( n3496 , n3423 , n3432 );
and ( n3497 , n3496 , n2899 );
or ( n3498 , n3495 , n3497 );
not ( n3499 , n3498 );
not ( n3500 , n3499 );
not ( n3501 , n3500 );
not ( n3502 , n2899 );
and ( n3503 , n3502 , n2779 );
xor ( n3504 , n3424 , n3431 );
and ( n3505 , n3504 , n2899 );
or ( n3506 , n3503 , n3505 );
not ( n3507 , n3506 );
not ( n3508 , n3507 );
not ( n3509 , n3508 );
not ( n3510 , n2899 );
and ( n3511 , n3510 , n2764 );
xor ( n3512 , n3425 , n3430 );
and ( n3513 , n3512 , n2899 );
or ( n3514 , n3511 , n3513 );
not ( n3515 , n3514 );
not ( n3516 , n3515 );
not ( n3517 , n3516 );
not ( n3518 , n2899 );
and ( n3519 , n3518 , n2749 );
xor ( n3520 , n3426 , n3429 );
and ( n3521 , n3520 , n2899 );
or ( n3522 , n3519 , n3521 );
not ( n3523 , n3522 );
not ( n3524 , n3523 );
not ( n3525 , n3524 );
not ( n3526 , n2899 );
and ( n3527 , n3526 , n2734 );
xor ( n3528 , n3427 , n3428 );
and ( n3529 , n3528 , n2899 );
or ( n3530 , n3527 , n3529 );
not ( n3531 , n3530 );
not ( n3532 , n3531 );
not ( n3533 , n3532 );
not ( n3534 , n3408 );
and ( n3535 , n3533 , n3534 );
and ( n3536 , n3525 , n3535 );
and ( n3537 , n3517 , n3536 );
and ( n3538 , n3509 , n3537 );
and ( n3539 , n3501 , n3538 );
and ( n3540 , n3493 , n3539 );
and ( n3541 , n3485 , n3540 );
and ( n3542 , n3477 , n3541 );
and ( n3543 , n3469 , n3542 );
and ( n3544 , n3461 , n3543 );
and ( n3545 , n3453 , n3544 );
and ( n3546 , n3445 , n3545 );
not ( n3547 , n3546 );
and ( n3548 , n3547 , n2899 );
or ( n3549 , n3412 , n3548 );
not ( n3550 , n3549 );
not ( n3551 , n2899 );
and ( n3552 , n3551 , n3532 );
xor ( n3553 , n3533 , n3534 );
and ( n3554 , n3553 , n2899 );
or ( n3555 , n3552 , n3554 );
and ( n3556 , n3550 , n3555 );
not ( n3557 , n3555 );
not ( n3558 , n3408 );
xor ( n3559 , n3557 , n3558 );
and ( n3560 , n3559 , n3549 );
or ( n3561 , n3556 , n3560 );
not ( n3562 , n3561 );
not ( n3563 , n3562 );
or ( n3564 , n3410 , n3563 );
not ( n3565 , n3549 );
not ( n3566 , n2899 );
and ( n3567 , n3566 , n3524 );
xor ( n3568 , n3525 , n3535 );
and ( n3569 , n3568 , n2899 );
or ( n3570 , n3567 , n3569 );
and ( n3571 , n3565 , n3570 );
not ( n3572 , n3570 );
and ( n3573 , n3557 , n3558 );
xor ( n3574 , n3572 , n3573 );
and ( n3575 , n3574 , n3549 );
or ( n3576 , n3571 , n3575 );
not ( n3577 , n3576 );
not ( n3578 , n3577 );
or ( n3579 , n3564 , n3578 );
not ( n3580 , n3549 );
not ( n3581 , n2899 );
and ( n3582 , n3581 , n3516 );
xor ( n3583 , n3517 , n3536 );
and ( n3584 , n3583 , n2899 );
or ( n3585 , n3582 , n3584 );
and ( n3586 , n3580 , n3585 );
not ( n3587 , n3585 );
and ( n3588 , n3572 , n3573 );
xor ( n3589 , n3587 , n3588 );
and ( n3590 , n3589 , n3549 );
or ( n3591 , n3586 , n3590 );
not ( n3592 , n3591 );
not ( n3593 , n3592 );
or ( n3594 , n3579 , n3593 );
buf ( n3595 , n3594 );
buf ( n3596 , n3595 );
and ( n3597 , n3596 , n3549 );
not ( n3598 , n3597 );
and ( n3599 , n3598 , n3410 );
xor ( n3600 , n3410 , n3549 );
xor ( n3601 , n3600 , n3549 );
and ( n3602 , n3601 , n3597 );
or ( n3603 , n3599 , n3602 );
not ( n3604 , n3597 );
and ( n3605 , n3604 , n3563 );
xor ( n3606 , n3563 , n3549 );
and ( n3607 , n3600 , n3549 );
xor ( n3608 , n3606 , n3607 );
and ( n3609 , n3608 , n3597 );
or ( n3610 , n3605 , n3609 );
not ( n3611 , n3610 );
not ( n3612 , n3597 );
and ( n3613 , n3612 , n3578 );
xor ( n3614 , n3578 , n3549 );
and ( n3615 , n3606 , n3607 );
xor ( n3616 , n3614 , n3615 );
and ( n3617 , n3616 , n3597 );
or ( n3618 , n3613 , n3617 );
not ( n3619 , n3597 );
and ( n3620 , n3619 , n3593 );
xor ( n3621 , n3593 , n3549 );
and ( n3622 , n3614 , n3615 );
xor ( n3623 , n3621 , n3622 );
and ( n3624 , n3623 , n3597 );
or ( n3625 , n3620 , n3624 );
and ( n3626 , n3603 , n3611 , n3618 , n3625 );
not ( n3627 , n3603 );
and ( n3628 , n3627 , n3610 , n3618 , n3625 );
or ( n3629 , n3626 , n3628 );
and ( n3630 , n3603 , n3610 , n3618 , n3625 );
or ( n3631 , n3629 , n3630 );
and ( n3632 , n3363 , n3631 );
buf ( n3633 , n2424 );
not ( n3634 , n3290 );
buf ( n3635 , n190 );
not ( n3636 , n2899 );
and ( n3637 , n3636 , n2869 );
not ( n3638 , n2869 );
not ( n3639 , n2854 );
not ( n3640 , n2839 );
not ( n3641 , n2824 );
not ( n3642 , n2809 );
not ( n3643 , n2794 );
not ( n3644 , n2779 );
not ( n3645 , n2764 );
not ( n3646 , n2749 );
not ( n3647 , n2734 );
not ( n3648 , n2719 );
not ( n3649 , n2704 );
not ( n3650 , n2689 );
not ( n3651 , n2674 );
not ( n3652 , n2659 );
not ( n3653 , n2644 );
not ( n3654 , n2629 );
not ( n3655 , n2614 );
not ( n3656 , n2599 );
not ( n3657 , n2584 );
not ( n3658 , n2569 );
not ( n3659 , n2554 );
not ( n3660 , n2539 );
not ( n3661 , n2524 );
not ( n3662 , n2509 );
not ( n3663 , n2494 );
not ( n3664 , n2479 );
not ( n3665 , n2464 );
not ( n3666 , n2449 );
not ( n3667 , n2430 );
and ( n3668 , n3666 , n3667 );
and ( n3669 , n3665 , n3668 );
and ( n3670 , n3664 , n3669 );
and ( n3671 , n3663 , n3670 );
and ( n3672 , n3662 , n3671 );
and ( n3673 , n3661 , n3672 );
and ( n3674 , n3660 , n3673 );
and ( n3675 , n3659 , n3674 );
and ( n3676 , n3658 , n3675 );
and ( n3677 , n3657 , n3676 );
and ( n3678 , n3656 , n3677 );
and ( n3679 , n3655 , n3678 );
and ( n3680 , n3654 , n3679 );
and ( n3681 , n3653 , n3680 );
and ( n3682 , n3652 , n3681 );
and ( n3683 , n3651 , n3682 );
and ( n3684 , n3650 , n3683 );
and ( n3685 , n3649 , n3684 );
and ( n3686 , n3648 , n3685 );
and ( n3687 , n3647 , n3686 );
and ( n3688 , n3646 , n3687 );
and ( n3689 , n3645 , n3688 );
and ( n3690 , n3644 , n3689 );
and ( n3691 , n3643 , n3690 );
and ( n3692 , n3642 , n3691 );
and ( n3693 , n3641 , n3692 );
and ( n3694 , n3640 , n3693 );
and ( n3695 , n3639 , n3694 );
xor ( n3696 , n3638 , n3695 );
and ( n3697 , n3696 , n2899 );
or ( n3698 , n3637 , n3697 );
not ( n3699 , n3698 );
not ( n3700 , n3699 );
not ( n3701 , n3700 );
not ( n3702 , n3701 );
not ( n3703 , n2899 );
and ( n3704 , n3703 , n2424 );
buf ( n3705 , n2899 );
not ( n3706 , n3705 );
and ( n3707 , n3706 , n2899 );
not ( n3708 , n2899 );
not ( n3709 , n2884 );
and ( n3710 , n3638 , n3695 );
and ( n3711 , n3709 , n3710 );
xor ( n3712 , n3708 , n3711 );
and ( n3713 , n3712 , n3705 );
or ( n3714 , n3707 , n3713 );
not ( n3715 , n3714 );
not ( n3716 , n3715 );
not ( n3717 , n3716 );
not ( n3718 , n2899 );
and ( n3719 , n3718 , n2884 );
xor ( n3720 , n3709 , n3710 );
and ( n3721 , n3720 , n2899 );
or ( n3722 , n3719 , n3721 );
not ( n3723 , n3722 );
not ( n3724 , n3723 );
not ( n3725 , n3724 );
not ( n3726 , n3700 );
and ( n3727 , n3725 , n3726 );
and ( n3728 , n3717 , n3727 );
not ( n3729 , n3728 );
and ( n3730 , n3729 , n2899 );
or ( n3731 , n3704 , n3730 );
not ( n3732 , n3731 );
not ( n3733 , n2899 );
and ( n3734 , n3733 , n3724 );
xor ( n3735 , n3725 , n3726 );
and ( n3736 , n3735 , n2899 );
or ( n3737 , n3734 , n3736 );
and ( n3738 , n3732 , n3737 );
not ( n3739 , n3737 );
not ( n3740 , n3700 );
xor ( n3741 , n3739 , n3740 );
and ( n3742 , n3741 , n3731 );
or ( n3743 , n3738 , n3742 );
not ( n3744 , n3743 );
not ( n3745 , n3744 );
or ( n3746 , n3702 , n3745 );
and ( n3747 , n3746 , n3731 );
not ( n3748 , n3747 );
and ( n3749 , n3748 , n3702 );
xor ( n3750 , n3702 , n3731 );
xor ( n3751 , n3750 , n3731 );
and ( n3752 , n3751 , n3747 );
or ( n3753 , n3749 , n3752 );
not ( n3754 , n3753 );
not ( n3755 , n3747 );
and ( n3756 , n3755 , n3745 );
xor ( n3757 , n3745 , n3731 );
and ( n3758 , n3750 , n3731 );
xor ( n3759 , n3757 , n3758 );
and ( n3760 , n3759 , n3747 );
or ( n3761 , n3756 , n3760 );
and ( n3762 , n3754 , n3761 );
and ( n3763 , n3635 , n3762 );
buf ( n3764 , n126 );
nor ( n3765 , n3754 , n3761 );
and ( n3766 , n3764 , n3765 );
buf ( n3767 , n158 );
nor ( n3768 , n3753 , n3761 );
and ( n3769 , n3767 , n3768 );
or ( n3770 , n2424 , n3763 , n3766 , n3769 );
not ( n3771 , n3770 );
buf ( n3772 , n67 );
buf ( n3773 , n3772 );
not ( n3774 , n3773 );
not ( n3775 , n3774 );
buf ( n3776 , n3775 );
and ( n3777 , n3753 , n3761 );
and ( n3778 , n3776 , n3777 );
buf ( n3779 , n160 );
and ( n3780 , n3779 , n3762 );
buf ( n3781 , n96 );
and ( n3782 , n3781 , n3765 );
buf ( n3783 , n128 );
and ( n3784 , n3783 , n3768 );
or ( n3785 , n3778 , n3780 , n3782 , n3784 );
and ( n3786 , n3771 , n3785 );
not ( n3787 , n3785 );
and ( n3788 , n3363 , n3777 );
buf ( n3789 , n159 );
and ( n3790 , n3789 , n3762 );
buf ( n3791 , n95 );
and ( n3792 , n3791 , n3765 );
buf ( n3793 , n127 );
and ( n3794 , n3793 , n3768 );
or ( n3795 , n3788 , n3790 , n3792 , n3794 );
not ( n3796 , n3795 );
xor ( n3797 , n3787 , n3796 );
and ( n3798 , n3797 , n3770 );
or ( n3799 , n3786 , n3798 );
not ( n3800 , n3799 );
buf ( n3801 , n3800 );
buf ( n3802 , n3801 );
not ( n3803 , n3802 );
and ( n3804 , n3634 , n3803 );
not ( n3805 , n3803 );
not ( n3806 , n3805 );
not ( n3807 , n3770 );
and ( n3808 , n3807 , n2424 );
buf ( n3809 , n3770 );
not ( n3810 , n3809 );
and ( n3811 , n3810 , n3770 );
not ( n3812 , n3770 );
buf ( n3813 , n189 );
and ( n3814 , n3813 , n3762 );
buf ( n3815 , n125 );
and ( n3816 , n3815 , n3765 );
buf ( n3817 , n157 );
and ( n3818 , n3817 , n3768 );
or ( n3819 , n2424 , n3814 , n3816 , n3818 );
not ( n3820 , n3819 );
buf ( n3821 , n94 );
buf ( n3822 , n3821 );
not ( n3823 , n3822 );
not ( n3824 , n3823 );
buf ( n3825 , n3824 );
buf ( n3826 , n93 );
buf ( n3827 , n3826 );
not ( n3828 , n3827 );
not ( n3829 , n3828 );
buf ( n3830 , n3829 );
buf ( n3831 , n92 );
buf ( n3832 , n3831 );
not ( n3833 , n3832 );
not ( n3834 , n3833 );
buf ( n3835 , n3834 );
buf ( n3836 , n91 );
buf ( n3837 , n3836 );
not ( n3838 , n3837 );
not ( n3839 , n3838 );
buf ( n3840 , n3839 );
buf ( n3841 , n90 );
buf ( n3842 , n3841 );
not ( n3843 , n3842 );
not ( n3844 , n3843 );
buf ( n3845 , n3844 );
buf ( n3846 , n89 );
buf ( n3847 , n3846 );
not ( n3848 , n3847 );
not ( n3849 , n3848 );
buf ( n3850 , n3849 );
buf ( n3851 , n88 );
buf ( n3852 , n3851 );
not ( n3853 , n3852 );
not ( n3854 , n3853 );
buf ( n3855 , n3854 );
buf ( n3856 , n87 );
buf ( n3857 , n3856 );
not ( n3858 , n3857 );
buf ( n3859 , n3858 );
buf ( n3860 , n86 );
buf ( n3861 , n3860 );
not ( n3862 , n3861 );
not ( n3863 , n3862 );
buf ( n3864 , n3863 );
buf ( n3865 , n85 );
buf ( n3866 , n3865 );
not ( n3867 , n3866 );
not ( n3868 , n3867 );
buf ( n3869 , n3868 );
buf ( n3870 , n84 );
buf ( n3871 , n3870 );
not ( n3872 , n3871 );
not ( n3873 , n3872 );
buf ( n3874 , n3873 );
buf ( n3875 , n83 );
buf ( n3876 , n3875 );
not ( n3877 , n3876 );
not ( n3878 , n3877 );
buf ( n3879 , n3878 );
buf ( n3880 , n82 );
buf ( n3881 , n3880 );
not ( n3882 , n3881 );
not ( n3883 , n3882 );
buf ( n3884 , n3883 );
buf ( n3885 , n81 );
buf ( n3886 , n3885 );
not ( n3887 , n3886 );
not ( n3888 , n3887 );
buf ( n3889 , n3888 );
buf ( n3890 , n80 );
buf ( n3891 , n3890 );
not ( n3892 , n3891 );
not ( n3893 , n3892 );
buf ( n3894 , n3893 );
buf ( n3895 , n79 );
buf ( n3896 , n3895 );
not ( n3897 , n3896 );
not ( n3898 , n3897 );
buf ( n3899 , n3898 );
buf ( n3900 , n78 );
buf ( n3901 , n3900 );
not ( n3902 , n3901 );
not ( n3903 , n3902 );
buf ( n3904 , n3903 );
buf ( n3905 , n77 );
buf ( n3906 , n3905 );
not ( n3907 , n3906 );
not ( n3908 , n3907 );
buf ( n3909 , n3908 );
buf ( n3910 , n76 );
buf ( n3911 , n3910 );
not ( n3912 , n3911 );
not ( n3913 , n3912 );
buf ( n3914 , n3913 );
buf ( n3915 , n75 );
buf ( n3916 , n3915 );
not ( n3917 , n3916 );
not ( n3918 , n3917 );
buf ( n3919 , n3918 );
buf ( n3920 , n74 );
buf ( n3921 , n3920 );
not ( n3922 , n3921 );
not ( n3923 , n3922 );
buf ( n3924 , n3923 );
buf ( n3925 , n73 );
buf ( n3926 , n3925 );
not ( n3927 , n3926 );
not ( n3928 , n3927 );
buf ( n3929 , n3928 );
buf ( n3930 , n72 );
buf ( n3931 , n3930 );
not ( n3932 , n3931 );
not ( n3933 , n3932 );
buf ( n3934 , n3933 );
buf ( n3935 , n71 );
buf ( n3936 , n3935 );
not ( n3937 , n3936 );
not ( n3938 , n3937 );
buf ( n3939 , n3938 );
buf ( n3940 , n70 );
buf ( n3941 , n3940 );
not ( n3942 , n3941 );
not ( n3943 , n3942 );
buf ( n3944 , n3943 );
buf ( n3945 , n69 );
buf ( n3946 , n3945 );
not ( n3947 , n3946 );
not ( n3948 , n3947 );
buf ( n3949 , n3948 );
and ( n3950 , n3944 , n3949 );
and ( n3951 , n3939 , n3950 );
and ( n3952 , n3934 , n3951 );
and ( n3953 , n3929 , n3952 );
and ( n3954 , n3924 , n3953 );
and ( n3955 , n3919 , n3954 );
and ( n3956 , n3914 , n3955 );
and ( n3957 , n3909 , n3956 );
and ( n3958 , n3904 , n3957 );
and ( n3959 , n3899 , n3958 );
and ( n3960 , n3894 , n3959 );
and ( n3961 , n3889 , n3960 );
and ( n3962 , n3884 , n3961 );
and ( n3963 , n3879 , n3962 );
and ( n3964 , n3874 , n3963 );
and ( n3965 , n3869 , n3964 );
and ( n3966 , n3864 , n3965 );
and ( n3967 , n3859 , n3966 );
and ( n3968 , n3855 , n3967 );
and ( n3969 , n3850 , n3968 );
and ( n3970 , n3845 , n3969 );
and ( n3971 , n3840 , n3970 );
and ( n3972 , n3835 , n3971 );
and ( n3973 , n3830 , n3972 );
and ( n3974 , n3825 , n3973 );
buf ( n3975 , n3974 );
and ( n3976 , n3975 , n3777 );
buf ( n3977 , n188 );
and ( n3978 , n3977 , n3762 );
buf ( n3979 , n124 );
and ( n3980 , n3979 , n3765 );
buf ( n3981 , n156 );
and ( n3982 , n3981 , n3768 );
or ( n3983 , n3976 , n3978 , n3980 , n3982 );
not ( n3984 , n3983 );
xor ( n3985 , n3825 , n3973 );
and ( n3986 , n3985 , n3777 );
buf ( n3987 , n187 );
and ( n3988 , n3987 , n3762 );
buf ( n3989 , n123 );
and ( n3990 , n3989 , n3765 );
buf ( n3991 , n155 );
and ( n3992 , n3991 , n3768 );
or ( n3993 , n3986 , n3988 , n3990 , n3992 );
not ( n3994 , n3993 );
xor ( n3995 , n3830 , n3972 );
and ( n3996 , n3995 , n3777 );
buf ( n3997 , n186 );
and ( n3998 , n3997 , n3762 );
buf ( n3999 , n122 );
and ( n4000 , n3999 , n3765 );
buf ( n4001 , n154 );
and ( n4002 , n4001 , n3768 );
or ( n4003 , n3996 , n3998 , n4000 , n4002 );
not ( n4004 , n4003 );
xor ( n4005 , n3835 , n3971 );
and ( n4006 , n4005 , n3777 );
buf ( n4007 , n185 );
and ( n4008 , n4007 , n3762 );
buf ( n4009 , n121 );
and ( n4010 , n4009 , n3765 );
buf ( n4011 , n153 );
and ( n4012 , n4011 , n3768 );
or ( n4013 , n4006 , n4008 , n4010 , n4012 );
not ( n4014 , n4013 );
xor ( n4015 , n3840 , n3970 );
and ( n4016 , n4015 , n3777 );
buf ( n4017 , n184 );
and ( n4018 , n4017 , n3762 );
buf ( n4019 , n120 );
and ( n4020 , n4019 , n3765 );
buf ( n4021 , n152 );
and ( n4022 , n4021 , n3768 );
or ( n4023 , n4016 , n4018 , n4020 , n4022 );
not ( n4024 , n4023 );
xor ( n4025 , n3845 , n3969 );
and ( n4026 , n4025 , n3777 );
buf ( n4027 , n183 );
and ( n4028 , n4027 , n3762 );
buf ( n4029 , n119 );
and ( n4030 , n4029 , n3765 );
buf ( n4031 , n151 );
and ( n4032 , n4031 , n3768 );
or ( n4033 , n4026 , n4028 , n4030 , n4032 );
not ( n4034 , n4033 );
xor ( n4035 , n3850 , n3968 );
and ( n4036 , n4035 , n3777 );
buf ( n4037 , n182 );
and ( n4038 , n4037 , n3762 );
buf ( n4039 , n118 );
and ( n4040 , n4039 , n3765 );
buf ( n4041 , n150 );
and ( n4042 , n4041 , n3768 );
or ( n4043 , n4036 , n4038 , n4040 , n4042 );
not ( n4044 , n4043 );
xor ( n4045 , n3855 , n3967 );
and ( n4046 , n4045 , n3777 );
buf ( n4047 , n181 );
and ( n4048 , n4047 , n3762 );
buf ( n4049 , n117 );
and ( n4050 , n4049 , n3765 );
buf ( n4051 , n149 );
and ( n4052 , n4051 , n3768 );
or ( n4053 , n4046 , n4048 , n4050 , n4052 );
not ( n4054 , n4053 );
xor ( n4055 , n3859 , n3966 );
and ( n4056 , n4055 , n3777 );
buf ( n4057 , n180 );
and ( n4058 , n4057 , n3762 );
buf ( n4059 , n116 );
and ( n4060 , n4059 , n3765 );
buf ( n4061 , n148 );
and ( n4062 , n4061 , n3768 );
or ( n4063 , n4056 , n4058 , n4060 , n4062 );
not ( n4064 , n4063 );
xor ( n4065 , n3864 , n3965 );
and ( n4066 , n4065 , n3777 );
buf ( n4067 , n179 );
and ( n4068 , n4067 , n3762 );
buf ( n4069 , n115 );
and ( n4070 , n4069 , n3765 );
buf ( n4071 , n147 );
and ( n4072 , n4071 , n3768 );
or ( n4073 , n4066 , n4068 , n4070 , n4072 );
not ( n4074 , n4073 );
xor ( n4075 , n3869 , n3964 );
and ( n4076 , n4075 , n3777 );
buf ( n4077 , n178 );
and ( n4078 , n4077 , n3762 );
buf ( n4079 , n114 );
and ( n4080 , n4079 , n3765 );
buf ( n4081 , n146 );
and ( n4082 , n4081 , n3768 );
or ( n4083 , n4076 , n4078 , n4080 , n4082 );
not ( n4084 , n4083 );
xor ( n4085 , n3874 , n3963 );
and ( n4086 , n4085 , n3777 );
buf ( n4087 , n177 );
and ( n4088 , n4087 , n3762 );
buf ( n4089 , n113 );
and ( n4090 , n4089 , n3765 );
buf ( n4091 , n145 );
and ( n4092 , n4091 , n3768 );
or ( n4093 , n4086 , n4088 , n4090 , n4092 );
not ( n4094 , n4093 );
xor ( n4095 , n3879 , n3962 );
and ( n4096 , n4095 , n3777 );
buf ( n4097 , n176 );
and ( n4098 , n4097 , n3762 );
buf ( n4099 , n112 );
and ( n4100 , n4099 , n3765 );
buf ( n4101 , n144 );
and ( n4102 , n4101 , n3768 );
or ( n4103 , n4096 , n4098 , n4100 , n4102 );
not ( n4104 , n4103 );
xor ( n4105 , n3884 , n3961 );
and ( n4106 , n4105 , n3777 );
buf ( n4107 , n175 );
and ( n4108 , n4107 , n3762 );
buf ( n4109 , n111 );
and ( n4110 , n4109 , n3765 );
buf ( n4111 , n143 );
and ( n4112 , n4111 , n3768 );
or ( n4113 , n4106 , n4108 , n4110 , n4112 );
not ( n4114 , n4113 );
xor ( n4115 , n3889 , n3960 );
and ( n4116 , n4115 , n3777 );
buf ( n4117 , n174 );
and ( n4118 , n4117 , n3762 );
buf ( n4119 , n110 );
and ( n4120 , n4119 , n3765 );
buf ( n4121 , n142 );
and ( n4122 , n4121 , n3768 );
or ( n4123 , n4116 , n4118 , n4120 , n4122 );
not ( n4124 , n4123 );
xor ( n4125 , n3894 , n3959 );
and ( n4126 , n4125 , n3777 );
buf ( n4127 , n173 );
and ( n4128 , n4127 , n3762 );
buf ( n4129 , n109 );
and ( n4130 , n4129 , n3765 );
buf ( n4131 , n141 );
and ( n4132 , n4131 , n3768 );
or ( n4133 , n4126 , n4128 , n4130 , n4132 );
not ( n4134 , n4133 );
xor ( n4135 , n3899 , n3958 );
and ( n4136 , n4135 , n3777 );
buf ( n4137 , n172 );
and ( n4138 , n4137 , n3762 );
buf ( n4139 , n108 );
and ( n4140 , n4139 , n3765 );
buf ( n4141 , n140 );
and ( n4142 , n4141 , n3768 );
or ( n4143 , n4136 , n4138 , n4140 , n4142 );
not ( n4144 , n4143 );
xor ( n4145 , n3904 , n3957 );
and ( n4146 , n4145 , n3777 );
buf ( n4147 , n171 );
and ( n4148 , n4147 , n3762 );
buf ( n4149 , n107 );
and ( n4150 , n4149 , n3765 );
buf ( n4151 , n139 );
and ( n4152 , n4151 , n3768 );
or ( n4153 , n4146 , n4148 , n4150 , n4152 );
not ( n4154 , n4153 );
xor ( n4155 , n3909 , n3956 );
and ( n4156 , n4155 , n3777 );
buf ( n4157 , n170 );
and ( n4158 , n4157 , n3762 );
buf ( n4159 , n106 );
and ( n4160 , n4159 , n3765 );
buf ( n4161 , n138 );
and ( n4162 , n4161 , n3768 );
or ( n4163 , n4156 , n4158 , n4160 , n4162 );
not ( n4164 , n4163 );
xor ( n4165 , n3914 , n3955 );
and ( n4166 , n4165 , n3777 );
buf ( n4167 , n169 );
and ( n4168 , n4167 , n3762 );
buf ( n4169 , n105 );
and ( n4170 , n4169 , n3765 );
buf ( n4171 , n137 );
and ( n4172 , n4171 , n3768 );
or ( n4173 , n4166 , n4168 , n4170 , n4172 );
not ( n4174 , n4173 );
xor ( n4175 , n3919 , n3954 );
and ( n4176 , n4175 , n3777 );
buf ( n4177 , n168 );
and ( n4178 , n4177 , n3762 );
buf ( n4179 , n104 );
and ( n4180 , n4179 , n3765 );
buf ( n4181 , n136 );
and ( n4182 , n4181 , n3768 );
or ( n4183 , n4176 , n4178 , n4180 , n4182 );
not ( n4184 , n4183 );
xor ( n4185 , n3924 , n3953 );
and ( n4186 , n4185 , n3777 );
buf ( n4187 , n167 );
and ( n4188 , n4187 , n3762 );
buf ( n4189 , n103 );
and ( n4190 , n4189 , n3765 );
buf ( n4191 , n135 );
and ( n4192 , n4191 , n3768 );
or ( n4193 , n4186 , n4188 , n4190 , n4192 );
not ( n4194 , n4193 );
xor ( n4195 , n3929 , n3952 );
and ( n4196 , n4195 , n3777 );
buf ( n4197 , n166 );
and ( n4198 , n4197 , n3762 );
buf ( n4199 , n102 );
and ( n4200 , n4199 , n3765 );
buf ( n4201 , n134 );
and ( n4202 , n4201 , n3768 );
or ( n4203 , n4196 , n4198 , n4200 , n4202 );
not ( n4204 , n4203 );
xor ( n4205 , n3934 , n3951 );
and ( n4206 , n4205 , n3777 );
buf ( n4207 , n165 );
and ( n4208 , n4207 , n3762 );
buf ( n4209 , n101 );
and ( n4210 , n4209 , n3765 );
buf ( n4211 , n133 );
and ( n4212 , n4211 , n3768 );
or ( n4213 , n4206 , n4208 , n4210 , n4212 );
not ( n4214 , n4213 );
xor ( n4215 , n3939 , n3950 );
and ( n4216 , n4215 , n3777 );
buf ( n4217 , n164 );
and ( n4218 , n4217 , n3762 );
buf ( n4219 , n100 );
and ( n4220 , n4219 , n3765 );
buf ( n4221 , n132 );
and ( n4222 , n4221 , n3768 );
or ( n4223 , n4216 , n4218 , n4220 , n4222 );
not ( n4224 , n4223 );
xor ( n4225 , n3944 , n3949 );
and ( n4226 , n4225 , n3777 );
buf ( n4227 , n163 );
and ( n4228 , n4227 , n3762 );
buf ( n4229 , n99 );
and ( n4230 , n4229 , n3765 );
buf ( n4231 , n131 );
and ( n4232 , n4231 , n3768 );
or ( n4233 , n4226 , n4228 , n4230 , n4232 );
not ( n4234 , n4233 );
not ( n4235 , n3949 );
and ( n4236 , n4235 , n3777 );
buf ( n4237 , n162 );
and ( n4238 , n4237 , n3762 );
buf ( n4239 , n98 );
and ( n4240 , n4239 , n3765 );
buf ( n4241 , n130 );
and ( n4242 , n4241 , n3768 );
or ( n4243 , n4236 , n4238 , n4240 , n4242 );
not ( n4244 , n4243 );
buf ( n4245 , n68 );
buf ( n4246 , n4245 );
not ( n4247 , n4246 );
not ( n4248 , n4247 );
buf ( n4249 , n4248 );
and ( n4250 , n4249 , n3777 );
buf ( n4251 , n161 );
and ( n4252 , n4251 , n3762 );
buf ( n4253 , n97 );
and ( n4254 , n4253 , n3765 );
buf ( n4255 , n129 );
and ( n4256 , n4255 , n3768 );
or ( n4257 , n4250 , n4252 , n4254 , n4256 );
not ( n4258 , n4257 );
and ( n4259 , n3787 , n3796 );
and ( n4260 , n4258 , n4259 );
and ( n4261 , n4244 , n4260 );
and ( n4262 , n4234 , n4261 );
and ( n4263 , n4224 , n4262 );
and ( n4264 , n4214 , n4263 );
and ( n4265 , n4204 , n4264 );
and ( n4266 , n4194 , n4265 );
and ( n4267 , n4184 , n4266 );
and ( n4268 , n4174 , n4267 );
and ( n4269 , n4164 , n4268 );
and ( n4270 , n4154 , n4269 );
and ( n4271 , n4144 , n4270 );
and ( n4272 , n4134 , n4271 );
and ( n4273 , n4124 , n4272 );
and ( n4274 , n4114 , n4273 );
and ( n4275 , n4104 , n4274 );
and ( n4276 , n4094 , n4275 );
and ( n4277 , n4084 , n4276 );
and ( n4278 , n4074 , n4277 );
and ( n4279 , n4064 , n4278 );
and ( n4280 , n4054 , n4279 );
and ( n4281 , n4044 , n4280 );
and ( n4282 , n4034 , n4281 );
and ( n4283 , n4024 , n4282 );
and ( n4284 , n4014 , n4283 );
and ( n4285 , n4004 , n4284 );
and ( n4286 , n3994 , n4285 );
and ( n4287 , n3984 , n4286 );
and ( n4288 , n3820 , n4287 );
xor ( n4289 , n3812 , n4288 );
and ( n4290 , n4289 , n3809 );
or ( n4291 , n3811 , n4290 );
not ( n4292 , n4291 );
not ( n4293 , n4292 );
not ( n4294 , n4293 );
not ( n4295 , n3770 );
and ( n4296 , n4295 , n3819 );
xor ( n4297 , n3820 , n4287 );
and ( n4298 , n4297 , n3770 );
or ( n4299 , n4296 , n4298 );
not ( n4300 , n4299 );
not ( n4301 , n4300 );
not ( n4302 , n4301 );
not ( n4303 , n3770 );
and ( n4304 , n4303 , n3983 );
xor ( n4305 , n3984 , n4286 );
and ( n4306 , n4305 , n3770 );
or ( n4307 , n4304 , n4306 );
not ( n4308 , n4307 );
not ( n4309 , n4308 );
not ( n4310 , n4309 );
not ( n4311 , n3770 );
and ( n4312 , n4311 , n3993 );
xor ( n4313 , n3994 , n4285 );
and ( n4314 , n4313 , n3770 );
or ( n4315 , n4312 , n4314 );
not ( n4316 , n4315 );
not ( n4317 , n4316 );
not ( n4318 , n4317 );
not ( n4319 , n3770 );
and ( n4320 , n4319 , n4003 );
xor ( n4321 , n4004 , n4284 );
and ( n4322 , n4321 , n3770 );
or ( n4323 , n4320 , n4322 );
not ( n4324 , n4323 );
not ( n4325 , n4324 );
not ( n4326 , n4325 );
not ( n4327 , n3770 );
and ( n4328 , n4327 , n4013 );
xor ( n4329 , n4014 , n4283 );
and ( n4330 , n4329 , n3770 );
or ( n4331 , n4328 , n4330 );
not ( n4332 , n4331 );
not ( n4333 , n4332 );
not ( n4334 , n4333 );
not ( n4335 , n3770 );
and ( n4336 , n4335 , n4023 );
xor ( n4337 , n4024 , n4282 );
and ( n4338 , n4337 , n3770 );
or ( n4339 , n4336 , n4338 );
not ( n4340 , n4339 );
not ( n4341 , n4340 );
not ( n4342 , n4341 );
not ( n4343 , n3770 );
and ( n4344 , n4343 , n4033 );
xor ( n4345 , n4034 , n4281 );
and ( n4346 , n4345 , n3770 );
or ( n4347 , n4344 , n4346 );
not ( n4348 , n4347 );
not ( n4349 , n4348 );
not ( n4350 , n4349 );
not ( n4351 , n3770 );
and ( n4352 , n4351 , n4043 );
xor ( n4353 , n4044 , n4280 );
and ( n4354 , n4353 , n3770 );
or ( n4355 , n4352 , n4354 );
not ( n4356 , n4355 );
not ( n4357 , n4356 );
not ( n4358 , n4357 );
not ( n4359 , n3770 );
and ( n4360 , n4359 , n4053 );
xor ( n4361 , n4054 , n4279 );
and ( n4362 , n4361 , n3770 );
or ( n4363 , n4360 , n4362 );
not ( n4364 , n4363 );
not ( n4365 , n4364 );
not ( n4366 , n4365 );
not ( n4367 , n3770 );
and ( n4368 , n4367 , n4063 );
xor ( n4369 , n4064 , n4278 );
and ( n4370 , n4369 , n3770 );
or ( n4371 , n4368 , n4370 );
not ( n4372 , n4371 );
not ( n4373 , n4372 );
not ( n4374 , n4373 );
not ( n4375 , n3770 );
and ( n4376 , n4375 , n4073 );
xor ( n4377 , n4074 , n4277 );
and ( n4378 , n4377 , n3770 );
or ( n4379 , n4376 , n4378 );
not ( n4380 , n4379 );
not ( n4381 , n4380 );
not ( n4382 , n4381 );
not ( n4383 , n3770 );
and ( n4384 , n4383 , n4083 );
xor ( n4385 , n4084 , n4276 );
and ( n4386 , n4385 , n3770 );
or ( n4387 , n4384 , n4386 );
not ( n4388 , n4387 );
not ( n4389 , n4388 );
not ( n4390 , n4389 );
not ( n4391 , n3770 );
and ( n4392 , n4391 , n4093 );
xor ( n4393 , n4094 , n4275 );
and ( n4394 , n4393 , n3770 );
or ( n4395 , n4392 , n4394 );
not ( n4396 , n4395 );
not ( n4397 , n4396 );
not ( n4398 , n4397 );
not ( n4399 , n3770 );
and ( n4400 , n4399 , n4103 );
xor ( n4401 , n4104 , n4274 );
and ( n4402 , n4401 , n3770 );
or ( n4403 , n4400 , n4402 );
not ( n4404 , n4403 );
not ( n4405 , n4404 );
not ( n4406 , n4405 );
not ( n4407 , n3770 );
and ( n4408 , n4407 , n4113 );
xor ( n4409 , n4114 , n4273 );
and ( n4410 , n4409 , n3770 );
or ( n4411 , n4408 , n4410 );
not ( n4412 , n4411 );
not ( n4413 , n4412 );
not ( n4414 , n4413 );
not ( n4415 , n3770 );
and ( n4416 , n4415 , n4123 );
xor ( n4417 , n4124 , n4272 );
and ( n4418 , n4417 , n3770 );
or ( n4419 , n4416 , n4418 );
not ( n4420 , n4419 );
not ( n4421 , n4420 );
not ( n4422 , n4421 );
not ( n4423 , n3770 );
and ( n4424 , n4423 , n4133 );
xor ( n4425 , n4134 , n4271 );
and ( n4426 , n4425 , n3770 );
or ( n4427 , n4424 , n4426 );
not ( n4428 , n4427 );
not ( n4429 , n4428 );
not ( n4430 , n4429 );
not ( n4431 , n3770 );
and ( n4432 , n4431 , n4143 );
xor ( n4433 , n4144 , n4270 );
and ( n4434 , n4433 , n3770 );
or ( n4435 , n4432 , n4434 );
not ( n4436 , n4435 );
not ( n4437 , n4436 );
not ( n4438 , n4437 );
not ( n4439 , n3770 );
and ( n4440 , n4439 , n4153 );
xor ( n4441 , n4154 , n4269 );
and ( n4442 , n4441 , n3770 );
or ( n4443 , n4440 , n4442 );
not ( n4444 , n4443 );
not ( n4445 , n4444 );
not ( n4446 , n4445 );
not ( n4447 , n3770 );
and ( n4448 , n4447 , n4163 );
xor ( n4449 , n4164 , n4268 );
and ( n4450 , n4449 , n3770 );
or ( n4451 , n4448 , n4450 );
not ( n4452 , n4451 );
not ( n4453 , n4452 );
not ( n4454 , n4453 );
not ( n4455 , n3770 );
and ( n4456 , n4455 , n4173 );
xor ( n4457 , n4174 , n4267 );
and ( n4458 , n4457 , n3770 );
or ( n4459 , n4456 , n4458 );
not ( n4460 , n4459 );
buf ( n4461 , n4460 );
buf ( n4462 , n4461 );
not ( n4463 , n4462 );
not ( n4464 , n4463 );
not ( n4465 , n3770 );
and ( n4466 , n4465 , n4183 );
xor ( n4467 , n4184 , n4266 );
and ( n4468 , n4467 , n3770 );
or ( n4469 , n4466 , n4468 );
not ( n4470 , n4469 );
buf ( n4471 , n4470 );
buf ( n4472 , n4471 );
not ( n4473 , n4472 );
not ( n4474 , n4473 );
not ( n4475 , n3770 );
and ( n4476 , n4475 , n4193 );
xor ( n4477 , n4194 , n4265 );
and ( n4478 , n4477 , n3770 );
or ( n4479 , n4476 , n4478 );
not ( n4480 , n4479 );
buf ( n4481 , n4480 );
buf ( n4482 , n4481 );
not ( n4483 , n4482 );
not ( n4484 , n4483 );
not ( n4485 , n3770 );
and ( n4486 , n4485 , n4203 );
xor ( n4487 , n4204 , n4264 );
and ( n4488 , n4487 , n3770 );
or ( n4489 , n4486 , n4488 );
not ( n4490 , n4489 );
buf ( n4491 , n4490 );
buf ( n4492 , n4491 );
not ( n4493 , n4492 );
not ( n4494 , n4493 );
not ( n4495 , n3770 );
and ( n4496 , n4495 , n4213 );
xor ( n4497 , n4214 , n4263 );
and ( n4498 , n4497 , n3770 );
or ( n4499 , n4496 , n4498 );
not ( n4500 , n4499 );
buf ( n4501 , n4500 );
buf ( n4502 , n4501 );
not ( n4503 , n4502 );
not ( n4504 , n4503 );
not ( n4505 , n3770 );
and ( n4506 , n4505 , n4223 );
xor ( n4507 , n4224 , n4262 );
and ( n4508 , n4507 , n3770 );
or ( n4509 , n4506 , n4508 );
not ( n4510 , n4509 );
buf ( n4511 , n4510 );
buf ( n4512 , n4511 );
not ( n4513 , n4512 );
not ( n4514 , n4513 );
not ( n4515 , n3770 );
and ( n4516 , n4515 , n4233 );
xor ( n4517 , n4234 , n4261 );
and ( n4518 , n4517 , n3770 );
or ( n4519 , n4516 , n4518 );
not ( n4520 , n4519 );
buf ( n4521 , n4520 );
buf ( n4522 , n4521 );
not ( n4523 , n4522 );
not ( n4524 , n4523 );
not ( n4525 , n3770 );
and ( n4526 , n4525 , n4243 );
xor ( n4527 , n4244 , n4260 );
and ( n4528 , n4527 , n3770 );
or ( n4529 , n4526 , n4528 );
not ( n4530 , n4529 );
buf ( n4531 , n4530 );
buf ( n4532 , n4531 );
not ( n4533 , n4532 );
not ( n4534 , n4533 );
not ( n4535 , n3770 );
and ( n4536 , n4535 , n4257 );
xor ( n4537 , n4258 , n4259 );
and ( n4538 , n4537 , n3770 );
or ( n4539 , n4536 , n4538 );
not ( n4540 , n4539 );
buf ( n4541 , n4540 );
buf ( n4542 , n4541 );
not ( n4543 , n4542 );
not ( n4544 , n4543 );
not ( n4545 , n3803 );
and ( n4546 , n4544 , n4545 );
and ( n4547 , n4534 , n4546 );
and ( n4548 , n4524 , n4547 );
and ( n4549 , n4514 , n4548 );
and ( n4550 , n4504 , n4549 );
and ( n4551 , n4494 , n4550 );
and ( n4552 , n4484 , n4551 );
and ( n4553 , n4474 , n4552 );
and ( n4554 , n4464 , n4553 );
and ( n4555 , n4454 , n4554 );
and ( n4556 , n4446 , n4555 );
and ( n4557 , n4438 , n4556 );
and ( n4558 , n4430 , n4557 );
and ( n4559 , n4422 , n4558 );
and ( n4560 , n4414 , n4559 );
and ( n4561 , n4406 , n4560 );
and ( n4562 , n4398 , n4561 );
and ( n4563 , n4390 , n4562 );
and ( n4564 , n4382 , n4563 );
and ( n4565 , n4374 , n4564 );
and ( n4566 , n4366 , n4565 );
and ( n4567 , n4358 , n4566 );
and ( n4568 , n4350 , n4567 );
and ( n4569 , n4342 , n4568 );
and ( n4570 , n4334 , n4569 );
and ( n4571 , n4326 , n4570 );
and ( n4572 , n4318 , n4571 );
and ( n4573 , n4310 , n4572 );
and ( n4574 , n4302 , n4573 );
and ( n4575 , n4294 , n4574 );
not ( n4576 , n4575 );
and ( n4577 , n4576 , n3770 );
or ( n4578 , n3808 , n4577 );
not ( n4579 , n4578 );
not ( n4580 , n3770 );
and ( n4581 , n4580 , n4543 );
xor ( n4582 , n4544 , n4545 );
and ( n4583 , n4582 , n3770 );
or ( n4584 , n4581 , n4583 );
and ( n4585 , n4579 , n4584 );
not ( n4586 , n4584 );
not ( n4587 , n3803 );
xor ( n4588 , n4586 , n4587 );
and ( n4589 , n4588 , n4578 );
or ( n4590 , n4585 , n4589 );
not ( n4591 , n4590 );
not ( n4592 , n4591 );
or ( n4593 , n3806 , n4592 );
not ( n4594 , n4578 );
not ( n4595 , n3770 );
and ( n4596 , n4595 , n4533 );
xor ( n4597 , n4534 , n4546 );
and ( n4598 , n4597 , n3770 );
or ( n4599 , n4596 , n4598 );
and ( n4600 , n4594 , n4599 );
not ( n4601 , n4599 );
and ( n4602 , n4586 , n4587 );
xor ( n4603 , n4601 , n4602 );
and ( n4604 , n4603 , n4578 );
or ( n4605 , n4600 , n4604 );
not ( n4606 , n4605 );
not ( n4607 , n4606 );
or ( n4608 , n4593 , n4607 );
not ( n4609 , n4578 );
not ( n4610 , n3770 );
and ( n4611 , n4610 , n4523 );
xor ( n4612 , n4524 , n4547 );
and ( n4613 , n4612 , n3770 );
or ( n4614 , n4611 , n4613 );
and ( n4615 , n4609 , n4614 );
not ( n4616 , n4614 );
and ( n4617 , n4601 , n4602 );
xor ( n4618 , n4616 , n4617 );
and ( n4619 , n4618 , n4578 );
or ( n4620 , n4615 , n4619 );
not ( n4621 , n4620 );
not ( n4622 , n4621 );
or ( n4623 , n4608 , n4622 );
not ( n4624 , n4578 );
not ( n4625 , n3770 );
and ( n4626 , n4625 , n4513 );
xor ( n4627 , n4514 , n4548 );
and ( n4628 , n4627 , n3770 );
or ( n4629 , n4626 , n4628 );
and ( n4630 , n4624 , n4629 );
not ( n4631 , n4629 );
and ( n4632 , n4616 , n4617 );
xor ( n4633 , n4631 , n4632 );
and ( n4634 , n4633 , n4578 );
or ( n4635 , n4630 , n4634 );
not ( n4636 , n4635 );
not ( n4637 , n4636 );
or ( n4638 , n4623 , n4637 );
not ( n4639 , n4578 );
not ( n4640 , n3770 );
and ( n4641 , n4640 , n4503 );
xor ( n4642 , n4504 , n4549 );
and ( n4643 , n4642 , n3770 );
or ( n4644 , n4641 , n4643 );
and ( n4645 , n4639 , n4644 );
not ( n4646 , n4644 );
and ( n4647 , n4631 , n4632 );
xor ( n4648 , n4646 , n4647 );
and ( n4649 , n4648 , n4578 );
or ( n4650 , n4645 , n4649 );
not ( n4651 , n4650 );
not ( n4652 , n4651 );
or ( n4653 , n4638 , n4652 );
not ( n4654 , n4578 );
not ( n4655 , n3770 );
and ( n4656 , n4655 , n4493 );
xor ( n4657 , n4494 , n4550 );
and ( n4658 , n4657 , n3770 );
or ( n4659 , n4656 , n4658 );
and ( n4660 , n4654 , n4659 );
not ( n4661 , n4659 );
and ( n4662 , n4646 , n4647 );
xor ( n4663 , n4661 , n4662 );
and ( n4664 , n4663 , n4578 );
or ( n4665 , n4660 , n4664 );
not ( n4666 , n4665 );
not ( n4667 , n4666 );
or ( n4668 , n4653 , n4667 );
not ( n4669 , n4578 );
not ( n4670 , n3770 );
and ( n4671 , n4670 , n4483 );
xor ( n4672 , n4484 , n4551 );
and ( n4673 , n4672 , n3770 );
or ( n4674 , n4671 , n4673 );
and ( n4675 , n4669 , n4674 );
not ( n4676 , n4674 );
and ( n4677 , n4661 , n4662 );
xor ( n4678 , n4676 , n4677 );
and ( n4679 , n4678 , n4578 );
or ( n4680 , n4675 , n4679 );
not ( n4681 , n4680 );
not ( n4682 , n4681 );
or ( n4683 , n4668 , n4682 );
not ( n4684 , n4578 );
not ( n4685 , n3770 );
and ( n4686 , n4685 , n4473 );
xor ( n4687 , n4474 , n4552 );
and ( n4688 , n4687 , n3770 );
or ( n4689 , n4686 , n4688 );
and ( n4690 , n4684 , n4689 );
not ( n4691 , n4689 );
and ( n4692 , n4676 , n4677 );
xor ( n4693 , n4691 , n4692 );
and ( n4694 , n4693 , n4578 );
or ( n4695 , n4690 , n4694 );
not ( n4696 , n4695 );
not ( n4697 , n4696 );
or ( n4698 , n4683 , n4697 );
not ( n4699 , n4578 );
not ( n4700 , n3770 );
and ( n4701 , n4700 , n4463 );
xor ( n4702 , n4464 , n4553 );
and ( n4703 , n4702 , n3770 );
or ( n4704 , n4701 , n4703 );
and ( n4705 , n4699 , n4704 );
not ( n4706 , n4704 );
and ( n4707 , n4691 , n4692 );
xor ( n4708 , n4706 , n4707 );
and ( n4709 , n4708 , n4578 );
or ( n4710 , n4705 , n4709 );
not ( n4711 , n4710 );
not ( n4712 , n4711 );
or ( n4713 , n4698 , n4712 );
not ( n4714 , n4578 );
not ( n4715 , n3770 );
and ( n4716 , n4715 , n4453 );
xor ( n4717 , n4454 , n4554 );
and ( n4718 , n4717 , n3770 );
or ( n4719 , n4716 , n4718 );
and ( n4720 , n4714 , n4719 );
not ( n4721 , n4719 );
and ( n4722 , n4706 , n4707 );
xor ( n4723 , n4721 , n4722 );
and ( n4724 , n4723 , n4578 );
or ( n4725 , n4720 , n4724 );
not ( n4726 , n4725 );
not ( n4727 , n4726 );
or ( n4728 , n4713 , n4727 );
not ( n4729 , n4578 );
not ( n4730 , n3770 );
and ( n4731 , n4730 , n4445 );
xor ( n4732 , n4446 , n4555 );
and ( n4733 , n4732 , n3770 );
or ( n4734 , n4731 , n4733 );
and ( n4735 , n4729 , n4734 );
not ( n4736 , n4734 );
and ( n4737 , n4721 , n4722 );
xor ( n4738 , n4736 , n4737 );
and ( n4739 , n4738 , n4578 );
or ( n4740 , n4735 , n4739 );
not ( n4741 , n4740 );
not ( n4742 , n4741 );
or ( n4743 , n4728 , n4742 );
not ( n4744 , n4578 );
not ( n4745 , n3770 );
and ( n4746 , n4745 , n4437 );
xor ( n4747 , n4438 , n4556 );
and ( n4748 , n4747 , n3770 );
or ( n4749 , n4746 , n4748 );
and ( n4750 , n4744 , n4749 );
not ( n4751 , n4749 );
and ( n4752 , n4736 , n4737 );
xor ( n4753 , n4751 , n4752 );
and ( n4754 , n4753 , n4578 );
or ( n4755 , n4750 , n4754 );
not ( n4756 , n4755 );
not ( n4757 , n4756 );
or ( n4758 , n4743 , n4757 );
not ( n4759 , n4578 );
not ( n4760 , n3770 );
and ( n4761 , n4760 , n4429 );
xor ( n4762 , n4430 , n4557 );
and ( n4763 , n4762 , n3770 );
or ( n4764 , n4761 , n4763 );
and ( n4765 , n4759 , n4764 );
not ( n4766 , n4764 );
and ( n4767 , n4751 , n4752 );
xor ( n4768 , n4766 , n4767 );
and ( n4769 , n4768 , n4578 );
or ( n4770 , n4765 , n4769 );
not ( n4771 , n4770 );
not ( n4772 , n4771 );
or ( n4773 , n4758 , n4772 );
not ( n4774 , n4578 );
not ( n4775 , n3770 );
and ( n4776 , n4775 , n4421 );
xor ( n4777 , n4422 , n4558 );
and ( n4778 , n4777 , n3770 );
or ( n4779 , n4776 , n4778 );
and ( n4780 , n4774 , n4779 );
not ( n4781 , n4779 );
and ( n4782 , n4766 , n4767 );
xor ( n4783 , n4781 , n4782 );
and ( n4784 , n4783 , n4578 );
or ( n4785 , n4780 , n4784 );
not ( n4786 , n4785 );
not ( n4787 , n4786 );
or ( n4788 , n4773 , n4787 );
not ( n4789 , n4578 );
not ( n4790 , n3770 );
and ( n4791 , n4790 , n4413 );
xor ( n4792 , n4414 , n4559 );
and ( n4793 , n4792 , n3770 );
or ( n4794 , n4791 , n4793 );
and ( n4795 , n4789 , n4794 );
not ( n4796 , n4794 );
and ( n4797 , n4781 , n4782 );
xor ( n4798 , n4796 , n4797 );
and ( n4799 , n4798 , n4578 );
or ( n4800 , n4795 , n4799 );
not ( n4801 , n4800 );
not ( n4802 , n4801 );
or ( n4803 , n4788 , n4802 );
not ( n4804 , n4578 );
not ( n4805 , n3770 );
and ( n4806 , n4805 , n4405 );
xor ( n4807 , n4406 , n4560 );
and ( n4808 , n4807 , n3770 );
or ( n4809 , n4806 , n4808 );
and ( n4810 , n4804 , n4809 );
not ( n4811 , n4809 );
and ( n4812 , n4796 , n4797 );
xor ( n4813 , n4811 , n4812 );
and ( n4814 , n4813 , n4578 );
or ( n4815 , n4810 , n4814 );
not ( n4816 , n4815 );
not ( n4817 , n4816 );
or ( n4818 , n4803 , n4817 );
not ( n4819 , n4578 );
not ( n4820 , n3770 );
and ( n4821 , n4820 , n4397 );
xor ( n4822 , n4398 , n4561 );
and ( n4823 , n4822 , n3770 );
or ( n4824 , n4821 , n4823 );
and ( n4825 , n4819 , n4824 );
not ( n4826 , n4824 );
and ( n4827 , n4811 , n4812 );
xor ( n4828 , n4826 , n4827 );
and ( n4829 , n4828 , n4578 );
or ( n4830 , n4825 , n4829 );
not ( n4831 , n4830 );
not ( n4832 , n4831 );
or ( n4833 , n4818 , n4832 );
not ( n4834 , n4578 );
not ( n4835 , n3770 );
and ( n4836 , n4835 , n4389 );
xor ( n4837 , n4390 , n4562 );
and ( n4838 , n4837 , n3770 );
or ( n4839 , n4836 , n4838 );
and ( n4840 , n4834 , n4839 );
not ( n4841 , n4839 );
and ( n4842 , n4826 , n4827 );
xor ( n4843 , n4841 , n4842 );
and ( n4844 , n4843 , n4578 );
or ( n4845 , n4840 , n4844 );
not ( n4846 , n4845 );
not ( n4847 , n4846 );
or ( n4848 , n4833 , n4847 );
not ( n4849 , n4578 );
not ( n4850 , n3770 );
and ( n4851 , n4850 , n4381 );
xor ( n4852 , n4382 , n4563 );
and ( n4853 , n4852 , n3770 );
or ( n4854 , n4851 , n4853 );
and ( n4855 , n4849 , n4854 );
not ( n4856 , n4854 );
and ( n4857 , n4841 , n4842 );
xor ( n4858 , n4856 , n4857 );
and ( n4859 , n4858 , n4578 );
or ( n4860 , n4855 , n4859 );
not ( n4861 , n4860 );
not ( n4862 , n4861 );
or ( n4863 , n4848 , n4862 );
not ( n4864 , n4578 );
not ( n4865 , n3770 );
and ( n4866 , n4865 , n4373 );
xor ( n4867 , n4374 , n4564 );
and ( n4868 , n4867 , n3770 );
or ( n4869 , n4866 , n4868 );
and ( n4870 , n4864 , n4869 );
not ( n4871 , n4869 );
and ( n4872 , n4856 , n4857 );
xor ( n4873 , n4871 , n4872 );
and ( n4874 , n4873 , n4578 );
or ( n4875 , n4870 , n4874 );
not ( n4876 , n4875 );
not ( n4877 , n4876 );
or ( n4878 , n4863 , n4877 );
not ( n4879 , n4578 );
not ( n4880 , n3770 );
and ( n4881 , n4880 , n4365 );
xor ( n4882 , n4366 , n4565 );
and ( n4883 , n4882 , n3770 );
or ( n4884 , n4881 , n4883 );
and ( n4885 , n4879 , n4884 );
not ( n4886 , n4884 );
and ( n4887 , n4871 , n4872 );
xor ( n4888 , n4886 , n4887 );
and ( n4889 , n4888 , n4578 );
or ( n4890 , n4885 , n4889 );
not ( n4891 , n4890 );
not ( n4892 , n4891 );
or ( n4893 , n4878 , n4892 );
not ( n4894 , n4578 );
not ( n4895 , n3770 );
and ( n4896 , n4895 , n4357 );
xor ( n4897 , n4358 , n4566 );
and ( n4898 , n4897 , n3770 );
or ( n4899 , n4896 , n4898 );
and ( n4900 , n4894 , n4899 );
not ( n4901 , n4899 );
and ( n4902 , n4886 , n4887 );
xor ( n4903 , n4901 , n4902 );
and ( n4904 , n4903 , n4578 );
or ( n4905 , n4900 , n4904 );
not ( n4906 , n4905 );
not ( n4907 , n4906 );
or ( n4908 , n4893 , n4907 );
not ( n4909 , n4578 );
not ( n4910 , n3770 );
and ( n4911 , n4910 , n4349 );
xor ( n4912 , n4350 , n4567 );
and ( n4913 , n4912 , n3770 );
or ( n4914 , n4911 , n4913 );
and ( n4915 , n4909 , n4914 );
not ( n4916 , n4914 );
and ( n4917 , n4901 , n4902 );
xor ( n4918 , n4916 , n4917 );
and ( n4919 , n4918 , n4578 );
or ( n4920 , n4915 , n4919 );
not ( n4921 , n4920 );
not ( n4922 , n4921 );
or ( n4923 , n4908 , n4922 );
not ( n4924 , n4578 );
not ( n4925 , n3770 );
and ( n4926 , n4925 , n4341 );
xor ( n4927 , n4342 , n4568 );
and ( n4928 , n4927 , n3770 );
or ( n4929 , n4926 , n4928 );
and ( n4930 , n4924 , n4929 );
not ( n4931 , n4929 );
and ( n4932 , n4916 , n4917 );
xor ( n4933 , n4931 , n4932 );
and ( n4934 , n4933 , n4578 );
or ( n4935 , n4930 , n4934 );
not ( n4936 , n4935 );
not ( n4937 , n4936 );
or ( n4938 , n4923 , n4937 );
not ( n4939 , n4578 );
not ( n4940 , n3770 );
and ( n4941 , n4940 , n4333 );
xor ( n4942 , n4334 , n4569 );
and ( n4943 , n4942 , n3770 );
or ( n4944 , n4941 , n4943 );
and ( n4945 , n4939 , n4944 );
not ( n4946 , n4944 );
and ( n4947 , n4931 , n4932 );
xor ( n4948 , n4946 , n4947 );
and ( n4949 , n4948 , n4578 );
or ( n4950 , n4945 , n4949 );
not ( n4951 , n4950 );
not ( n4952 , n4951 );
or ( n4953 , n4938 , n4952 );
not ( n4954 , n4578 );
not ( n4955 , n3770 );
and ( n4956 , n4955 , n4325 );
xor ( n4957 , n4326 , n4570 );
and ( n4958 , n4957 , n3770 );
or ( n4959 , n4956 , n4958 );
and ( n4960 , n4954 , n4959 );
not ( n4961 , n4959 );
and ( n4962 , n4946 , n4947 );
xor ( n4963 , n4961 , n4962 );
and ( n4964 , n4963 , n4578 );
or ( n4965 , n4960 , n4964 );
not ( n4966 , n4965 );
not ( n4967 , n4966 );
or ( n4968 , n4953 , n4967 );
not ( n4969 , n4578 );
not ( n4970 , n3770 );
and ( n4971 , n4970 , n4317 );
xor ( n4972 , n4318 , n4571 );
and ( n4973 , n4972 , n3770 );
or ( n4974 , n4971 , n4973 );
and ( n4975 , n4969 , n4974 );
not ( n4976 , n4974 );
and ( n4977 , n4961 , n4962 );
xor ( n4978 , n4976 , n4977 );
and ( n4979 , n4978 , n4578 );
or ( n4980 , n4975 , n4979 );
not ( n4981 , n4980 );
not ( n4982 , n4981 );
or ( n4983 , n4968 , n4982 );
not ( n4984 , n4578 );
not ( n4985 , n3770 );
and ( n4986 , n4985 , n4309 );
xor ( n4987 , n4310 , n4572 );
and ( n4988 , n4987 , n3770 );
or ( n4989 , n4986 , n4988 );
and ( n4990 , n4984 , n4989 );
not ( n4991 , n4989 );
and ( n4992 , n4976 , n4977 );
xor ( n4993 , n4991 , n4992 );
and ( n4994 , n4993 , n4578 );
or ( n4995 , n4990 , n4994 );
not ( n4996 , n4995 );
not ( n4997 , n4996 );
or ( n4998 , n4983 , n4997 );
and ( n4999 , n4998 , n4578 );
not ( n5000 , n4999 );
and ( n5001 , n5000 , n3806 );
xor ( n5002 , n3806 , n4578 );
xor ( n5003 , n5002 , n4578 );
and ( n5004 , n5003 , n4999 );
or ( n5005 , n5001 , n5004 );
and ( n5006 , n5005 , n3290 );
or ( n5007 , n3804 , n5006 );
not ( n5008 , n2899 );
and ( n5009 , n5008 , n2839 );
not ( n5010 , n2839 );
not ( n5011 , n2824 );
not ( n5012 , n2809 );
not ( n5013 , n2794 );
not ( n5014 , n2779 );
not ( n5015 , n2764 );
not ( n5016 , n2749 );
not ( n5017 , n2734 );
not ( n5018 , n2719 );
not ( n5019 , n2704 );
not ( n5020 , n2689 );
not ( n5021 , n2674 );
not ( n5022 , n2659 );
not ( n5023 , n2644 );
not ( n5024 , n2629 );
not ( n5025 , n2614 );
not ( n5026 , n2599 );
not ( n5027 , n2584 );
not ( n5028 , n2569 );
not ( n5029 , n2554 );
not ( n5030 , n2539 );
not ( n5031 , n2524 );
not ( n5032 , n2509 );
not ( n5033 , n2494 );
not ( n5034 , n2479 );
not ( n5035 , n2464 );
not ( n5036 , n2449 );
not ( n5037 , n2430 );
and ( n5038 , n5036 , n5037 );
and ( n5039 , n5035 , n5038 );
and ( n5040 , n5034 , n5039 );
and ( n5041 , n5033 , n5040 );
and ( n5042 , n5032 , n5041 );
and ( n5043 , n5031 , n5042 );
and ( n5044 , n5030 , n5043 );
and ( n5045 , n5029 , n5044 );
and ( n5046 , n5028 , n5045 );
and ( n5047 , n5027 , n5046 );
and ( n5048 , n5026 , n5047 );
and ( n5049 , n5025 , n5048 );
and ( n5050 , n5024 , n5049 );
and ( n5051 , n5023 , n5050 );
and ( n5052 , n5022 , n5051 );
and ( n5053 , n5021 , n5052 );
and ( n5054 , n5020 , n5053 );
and ( n5055 , n5019 , n5054 );
and ( n5056 , n5018 , n5055 );
and ( n5057 , n5017 , n5056 );
and ( n5058 , n5016 , n5057 );
and ( n5059 , n5015 , n5058 );
and ( n5060 , n5014 , n5059 );
and ( n5061 , n5013 , n5060 );
and ( n5062 , n5012 , n5061 );
and ( n5063 , n5011 , n5062 );
xor ( n5064 , n5010 , n5063 );
and ( n5065 , n5064 , n2899 );
or ( n5066 , n5009 , n5065 );
not ( n5067 , n5066 );
not ( n5068 , n5067 );
not ( n5069 , n5068 );
not ( n5070 , n5069 );
not ( n5071 , n2899 );
and ( n5072 , n5071 , n2424 );
buf ( n5073 , n2899 );
not ( n5074 , n5073 );
and ( n5075 , n5074 , n2899 );
not ( n5076 , n2899 );
not ( n5077 , n2884 );
not ( n5078 , n2869 );
not ( n5079 , n2854 );
and ( n5080 , n5010 , n5063 );
and ( n5081 , n5079 , n5080 );
and ( n5082 , n5078 , n5081 );
and ( n5083 , n5077 , n5082 );
xor ( n5084 , n5076 , n5083 );
and ( n5085 , n5084 , n5073 );
or ( n5086 , n5075 , n5085 );
not ( n5087 , n5086 );
not ( n5088 , n5087 );
not ( n5089 , n5088 );
not ( n5090 , n2899 );
and ( n5091 , n5090 , n2884 );
xor ( n5092 , n5077 , n5082 );
and ( n5093 , n5092 , n2899 );
or ( n5094 , n5091 , n5093 );
not ( n5095 , n5094 );
not ( n5096 , n5095 );
not ( n5097 , n5096 );
not ( n5098 , n2899 );
and ( n5099 , n5098 , n2869 );
xor ( n5100 , n5078 , n5081 );
and ( n5101 , n5100 , n2899 );
or ( n5102 , n5099 , n5101 );
not ( n5103 , n5102 );
not ( n5104 , n5103 );
not ( n5105 , n5104 );
not ( n5106 , n2899 );
and ( n5107 , n5106 , n2854 );
xor ( n5108 , n5079 , n5080 );
and ( n5109 , n5108 , n2899 );
or ( n5110 , n5107 , n5109 );
not ( n5111 , n5110 );
not ( n5112 , n5111 );
not ( n5113 , n5112 );
not ( n5114 , n5068 );
and ( n5115 , n5113 , n5114 );
and ( n5116 , n5105 , n5115 );
and ( n5117 , n5097 , n5116 );
and ( n5118 , n5089 , n5117 );
not ( n5119 , n5118 );
and ( n5120 , n5119 , n2899 );
or ( n5121 , n5072 , n5120 );
not ( n5122 , n5121 );
not ( n5123 , n2899 );
and ( n5124 , n5123 , n5112 );
xor ( n5125 , n5113 , n5114 );
and ( n5126 , n5125 , n2899 );
or ( n5127 , n5124 , n5126 );
and ( n5128 , n5122 , n5127 );
not ( n5129 , n5127 );
not ( n5130 , n5068 );
xor ( n5131 , n5129 , n5130 );
and ( n5132 , n5131 , n5121 );
or ( n5133 , n5128 , n5132 );
not ( n5134 , n5133 );
not ( n5135 , n5134 );
or ( n5136 , n5070 , n5135 );
and ( n5137 , n5136 , n5121 );
not ( n5138 , n5137 );
and ( n5139 , n5138 , n5070 );
xor ( n5140 , n5070 , n5121 );
xor ( n5141 , n5140 , n5121 );
and ( n5142 , n5141 , n5137 );
or ( n5143 , n5139 , n5142 );
not ( n5144 , n5143 );
not ( n5145 , n5137 );
and ( n5146 , n5145 , n5135 );
xor ( n5147 , n5135 , n5121 );
and ( n5148 , n5140 , n5121 );
xor ( n5149 , n5147 , n5148 );
and ( n5150 , n5149 , n5137 );
or ( n5151 , n5146 , n5150 );
nor ( n5152 , n5144 , n5151 );
and ( n5153 , n5007 , n5152 );
nor ( n5154 , n5143 , n5151 );
and ( n5155 , n3803 , n5154 );
or ( n5156 , n2424 , n3633 , n5153 , n5155 );
not ( n5157 , n3304 );
not ( n5158 , n3348 );
buf ( n5159 , n2424 );
buf ( n5160 , n2424 );
buf ( n5161 , n2424 );
buf ( n5162 , n2424 );
buf ( n5163 , n2424 );
buf ( n5164 , n2424 );
buf ( n5165 , n2424 );
buf ( n5166 , n2424 );
buf ( n5167 , n2424 );
buf ( n5168 , n2424 );
buf ( n5169 , n2424 );
buf ( n5170 , n2424 );
buf ( n5171 , n2424 );
buf ( n5172 , n2424 );
buf ( n5173 , n2424 );
buf ( n5174 , n2424 );
buf ( n5175 , n2424 );
buf ( n5176 , n2424 );
buf ( n5177 , n2424 );
buf ( n5178 , n2424 );
buf ( n5179 , n2424 );
buf ( n5180 , n2424 );
buf ( n5181 , n2424 );
buf ( n5182 , n2424 );
buf ( n5183 , n2424 );
buf ( n5184 , n2424 );
buf ( n5185 , n2424 );
buf ( n5186 , n2424 );
buf ( n5187 , n2424 );
nor ( n5188 , n5157 , n5158 , n2424 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 );
and ( n5189 , n5156 , n5188 );
buf ( n5190 , n2424 );
buf ( n5191 , n2424 );
buf ( n5192 , n2424 );
buf ( n5193 , n2424 );
buf ( n5194 , n2424 );
buf ( n5195 , n2424 );
buf ( n5196 , n2424 );
buf ( n5197 , n2424 );
buf ( n5198 , n2424 );
buf ( n5199 , n2424 );
buf ( n5200 , n2424 );
buf ( n5201 , n2424 );
buf ( n5202 , n2424 );
buf ( n5203 , n2424 );
buf ( n5204 , n2424 );
buf ( n5205 , n2424 );
buf ( n5206 , n2424 );
buf ( n5207 , n2424 );
buf ( n5208 , n2424 );
buf ( n5209 , n2424 );
buf ( n5210 , n2424 );
buf ( n5211 , n2424 );
buf ( n5212 , n2424 );
buf ( n5213 , n2424 );
buf ( n5214 , n2424 );
buf ( n5215 , n2424 );
buf ( n5216 , n2424 );
buf ( n5217 , n2424 );
buf ( n5218 , n2424 );
nor ( n5219 , n5157 , n3348 , n2424 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 );
buf ( n5220 , n2424 );
buf ( n5221 , n2424 );
buf ( n5222 , n2424 );
buf ( n5223 , n2424 );
buf ( n5224 , n2424 );
buf ( n5225 , n2424 );
buf ( n5226 , n2424 );
buf ( n5227 , n2424 );
buf ( n5228 , n2424 );
buf ( n5229 , n2424 );
buf ( n5230 , n2424 );
buf ( n5231 , n2424 );
buf ( n5232 , n2424 );
buf ( n5233 , n2424 );
buf ( n5234 , n2424 );
buf ( n5235 , n2424 );
buf ( n5236 , n2424 );
buf ( n5237 , n2424 );
buf ( n5238 , n2424 );
buf ( n5239 , n2424 );
buf ( n5240 , n2424 );
buf ( n5241 , n2424 );
buf ( n5242 , n2424 );
buf ( n5243 , n2424 );
buf ( n5244 , n2424 );
buf ( n5245 , n2424 );
buf ( n5246 , n2424 );
buf ( n5247 , n2424 );
buf ( n5248 , n2424 );
nor ( n5249 , n3304 , n3348 , n2424 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 );
or ( n5250 , n5219 , n5249 );
buf ( n5251 , n2424 );
buf ( n5252 , n2424 );
buf ( n5253 , n2424 );
buf ( n5254 , n2424 );
buf ( n5255 , n2424 );
buf ( n5256 , n2424 );
buf ( n5257 , n2424 );
buf ( n5258 , n2424 );
buf ( n5259 , n2424 );
buf ( n5260 , n2424 );
buf ( n5261 , n2424 );
buf ( n5262 , n2424 );
buf ( n5263 , n2424 );
buf ( n5264 , n2424 );
buf ( n5265 , n2424 );
buf ( n5266 , n2424 );
buf ( n5267 , n2424 );
buf ( n5268 , n2424 );
buf ( n5269 , n2424 );
buf ( n5270 , n2424 );
buf ( n5271 , n2424 );
buf ( n5272 , n2424 );
buf ( n5273 , n2424 );
buf ( n5274 , n2424 );
buf ( n5275 , n2424 );
buf ( n5276 , n2424 );
buf ( n5277 , n2424 );
buf ( n5278 , n2424 );
buf ( n5279 , n2424 );
nor ( n5280 , n3304 , n5158 , n2424 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 );
or ( n5281 , n5250 , n5280 );
buf ( n5282 , n5281 );
and ( n5283 , n3363 , n5282 );
or ( n5284 , n5189 , n5283 );
and ( n5285 , n3627 , n3611 , n3618 , n3625 );
and ( n5286 , n5284 , n5285 );
and ( n5287 , n5144 , n5151 );
or ( n5288 , n5152 , n5287 );
and ( n5289 , n5143 , n5151 );
or ( n5290 , n5288 , n5289 );
and ( n5291 , n2313 , n5290 );
not ( n5292 , n2430 );
not ( n5293 , n5292 );
not ( n5294 , n2899 );
and ( n5295 , n5294 , n2449 );
not ( n5296 , n2449 );
not ( n5297 , n2430 );
xor ( n5298 , n5296 , n5297 );
and ( n5299 , n5298 , n2899 );
or ( n5300 , n5295 , n5299 );
not ( n5301 , n5300 );
not ( n5302 , n5301 );
or ( n5303 , n5293 , n5302 );
not ( n5304 , n2899 );
and ( n5305 , n5304 , n2464 );
not ( n5306 , n2464 );
and ( n5307 , n5296 , n5297 );
xor ( n5308 , n5306 , n5307 );
and ( n5309 , n5308 , n2899 );
or ( n5310 , n5305 , n5309 );
not ( n5311 , n5310 );
not ( n5312 , n5311 );
or ( n5313 , n5303 , n5312 );
not ( n5314 , n2899 );
and ( n5315 , n5314 , n2479 );
not ( n5316 , n2479 );
and ( n5317 , n5306 , n5307 );
xor ( n5318 , n5316 , n5317 );
and ( n5319 , n5318 , n2899 );
or ( n5320 , n5315 , n5319 );
not ( n5321 , n5320 );
not ( n5322 , n5321 );
or ( n5323 , n5313 , n5322 );
not ( n5324 , n2899 );
and ( n5325 , n5324 , n2494 );
not ( n5326 , n2494 );
and ( n5327 , n5316 , n5317 );
xor ( n5328 , n5326 , n5327 );
and ( n5329 , n5328 , n2899 );
or ( n5330 , n5325 , n5329 );
not ( n5331 , n5330 );
not ( n5332 , n5331 );
or ( n5333 , n5323 , n5332 );
not ( n5334 , n2899 );
and ( n5335 , n5334 , n2509 );
not ( n5336 , n2509 );
and ( n5337 , n5326 , n5327 );
xor ( n5338 , n5336 , n5337 );
and ( n5339 , n5338 , n2899 );
or ( n5340 , n5335 , n5339 );
not ( n5341 , n5340 );
not ( n5342 , n5341 );
or ( n5343 , n5333 , n5342 );
not ( n5344 , n2899 );
and ( n5345 , n5344 , n2524 );
not ( n5346 , n2524 );
and ( n5347 , n5336 , n5337 );
xor ( n5348 , n5346 , n5347 );
and ( n5349 , n5348 , n2899 );
or ( n5350 , n5345 , n5349 );
not ( n5351 , n5350 );
not ( n5352 , n5351 );
or ( n5353 , n5343 , n5352 );
not ( n5354 , n2899 );
and ( n5355 , n5354 , n2539 );
not ( n5356 , n2539 );
and ( n5357 , n5346 , n5347 );
xor ( n5358 , n5356 , n5357 );
and ( n5359 , n5358 , n2899 );
or ( n5360 , n5355 , n5359 );
not ( n5361 , n5360 );
not ( n5362 , n5361 );
or ( n5363 , n5353 , n5362 );
not ( n5364 , n2899 );
and ( n5365 , n5364 , n2554 );
not ( n5366 , n2554 );
and ( n5367 , n5356 , n5357 );
xor ( n5368 , n5366 , n5367 );
and ( n5369 , n5368 , n2899 );
or ( n5370 , n5365 , n5369 );
not ( n5371 , n5370 );
not ( n5372 , n5371 );
or ( n5373 , n5363 , n5372 );
not ( n5374 , n2899 );
and ( n5375 , n5374 , n2569 );
not ( n5376 , n2569 );
and ( n5377 , n5366 , n5367 );
xor ( n5378 , n5376 , n5377 );
and ( n5379 , n5378 , n2899 );
or ( n5380 , n5375 , n5379 );
not ( n5381 , n5380 );
not ( n5382 , n5381 );
or ( n5383 , n5373 , n5382 );
not ( n5384 , n2899 );
and ( n5385 , n5384 , n2584 );
not ( n5386 , n2584 );
and ( n5387 , n5376 , n5377 );
xor ( n5388 , n5386 , n5387 );
and ( n5389 , n5388 , n2899 );
or ( n5390 , n5385 , n5389 );
not ( n5391 , n5390 );
not ( n5392 , n5391 );
or ( n5393 , n5383 , n5392 );
not ( n5394 , n2899 );
and ( n5395 , n5394 , n2599 );
not ( n5396 , n2599 );
and ( n5397 , n5386 , n5387 );
xor ( n5398 , n5396 , n5397 );
and ( n5399 , n5398 , n2899 );
or ( n5400 , n5395 , n5399 );
not ( n5401 , n5400 );
not ( n5402 , n5401 );
or ( n5403 , n5393 , n5402 );
not ( n5404 , n2899 );
and ( n5405 , n5404 , n2614 );
not ( n5406 , n2614 );
and ( n5407 , n5396 , n5397 );
xor ( n5408 , n5406 , n5407 );
and ( n5409 , n5408 , n2899 );
or ( n5410 , n5405 , n5409 );
not ( n5411 , n5410 );
not ( n5412 , n5411 );
or ( n5413 , n5403 , n5412 );
not ( n5414 , n2899 );
and ( n5415 , n5414 , n2629 );
not ( n5416 , n2629 );
and ( n5417 , n5406 , n5407 );
xor ( n5418 , n5416 , n5417 );
and ( n5419 , n5418 , n2899 );
or ( n5420 , n5415 , n5419 );
not ( n5421 , n5420 );
not ( n5422 , n5421 );
or ( n5423 , n5413 , n5422 );
not ( n5424 , n2899 );
and ( n5425 , n5424 , n2644 );
not ( n5426 , n2644 );
and ( n5427 , n5416 , n5417 );
xor ( n5428 , n5426 , n5427 );
and ( n5429 , n5428 , n2899 );
or ( n5430 , n5425 , n5429 );
not ( n5431 , n5430 );
not ( n5432 , n5431 );
or ( n5433 , n5423 , n5432 );
not ( n5434 , n2899 );
and ( n5435 , n5434 , n2659 );
not ( n5436 , n2659 );
and ( n5437 , n5426 , n5427 );
xor ( n5438 , n5436 , n5437 );
and ( n5439 , n5438 , n2899 );
or ( n5440 , n5435 , n5439 );
not ( n5441 , n5440 );
not ( n5442 , n5441 );
or ( n5443 , n5433 , n5442 );
not ( n5444 , n2899 );
and ( n5445 , n5444 , n2674 );
not ( n5446 , n2674 );
and ( n5447 , n5436 , n5437 );
xor ( n5448 , n5446 , n5447 );
and ( n5449 , n5448 , n2899 );
or ( n5450 , n5445 , n5449 );
not ( n5451 , n5450 );
not ( n5452 , n5451 );
or ( n5453 , n5443 , n5452 );
not ( n5454 , n2899 );
and ( n5455 , n5454 , n2689 );
not ( n5456 , n2689 );
and ( n5457 , n5446 , n5447 );
xor ( n5458 , n5456 , n5457 );
and ( n5459 , n5458 , n2899 );
or ( n5460 , n5455 , n5459 );
not ( n5461 , n5460 );
not ( n5462 , n5461 );
or ( n5463 , n5453 , n5462 );
not ( n5464 , n2899 );
and ( n5465 , n5464 , n2704 );
not ( n5466 , n2704 );
and ( n5467 , n5456 , n5457 );
xor ( n5468 , n5466 , n5467 );
and ( n5469 , n5468 , n2899 );
or ( n5470 , n5465 , n5469 );
not ( n5471 , n5470 );
not ( n5472 , n5471 );
or ( n5473 , n5463 , n5472 );
not ( n5474 , n2899 );
and ( n5475 , n5474 , n2719 );
not ( n5476 , n2719 );
and ( n5477 , n5466 , n5467 );
xor ( n5478 , n5476 , n5477 );
and ( n5479 , n5478 , n2899 );
or ( n5480 , n5475 , n5479 );
not ( n5481 , n5480 );
not ( n5482 , n5481 );
or ( n5483 , n5473 , n5482 );
and ( n5484 , n5483 , n2899 );
not ( n5485 , n5484 );
and ( n5486 , n5485 , n5293 );
xor ( n5487 , n5293 , n2899 );
xor ( n5488 , n5487 , n2899 );
and ( n5489 , n5488 , n5484 );
or ( n5490 , n5486 , n5489 );
and ( n5491 , n5490 , n5154 );
or ( n5492 , n5291 , n5491 );
xor ( n5493 , n3795 , n5492 );
not ( n5494 , n5493 );
not ( n5495 , n5494 );
and ( n5496 , n2282 , n5290 );
not ( n5497 , n5496 );
xor ( n5498 , n3770 , n5497 );
and ( n5499 , n2283 , n5290 );
not ( n5500 , n5499 );
and ( n5501 , n3819 , n5500 );
and ( n5502 , n2284 , n5290 );
not ( n5503 , n5502 );
and ( n5504 , n3983 , n5503 );
and ( n5505 , n2285 , n5290 );
not ( n5506 , n5505 );
and ( n5507 , n3993 , n5506 );
and ( n5508 , n2286 , n5290 );
not ( n5509 , n5508 );
and ( n5510 , n4003 , n5509 );
and ( n5511 , n2287 , n5290 );
not ( n5512 , n5511 );
and ( n5513 , n4013 , n5512 );
and ( n5514 , n2288 , n5290 );
not ( n5515 , n5514 );
and ( n5516 , n4023 , n5515 );
and ( n5517 , n2289 , n5290 );
not ( n5518 , n5517 );
and ( n5519 , n4033 , n5518 );
and ( n5520 , n2290 , n5290 );
not ( n5521 , n5520 );
and ( n5522 , n4043 , n5521 );
and ( n5523 , n2291 , n5290 );
not ( n5524 , n5523 );
and ( n5525 , n4053 , n5524 );
and ( n5526 , n2292 , n5290 );
not ( n5527 , n5526 );
and ( n5528 , n4063 , n5527 );
and ( n5529 , n2293 , n5290 );
not ( n5530 , n5529 );
and ( n5531 , n4073 , n5530 );
and ( n5532 , n2294 , n5290 );
not ( n5533 , n5484 );
and ( n5534 , n5533 , n5482 );
xor ( n5535 , n5482 , n2899 );
xor ( n5536 , n5472 , n2899 );
xor ( n5537 , n5462 , n2899 );
xor ( n5538 , n5452 , n2899 );
xor ( n5539 , n5442 , n2899 );
xor ( n5540 , n5432 , n2899 );
xor ( n5541 , n5422 , n2899 );
xor ( n5542 , n5412 , n2899 );
xor ( n5543 , n5402 , n2899 );
xor ( n5544 , n5392 , n2899 );
xor ( n5545 , n5382 , n2899 );
xor ( n5546 , n5372 , n2899 );
xor ( n5547 , n5362 , n2899 );
xor ( n5548 , n5352 , n2899 );
xor ( n5549 , n5342 , n2899 );
xor ( n5550 , n5332 , n2899 );
xor ( n5551 , n5322 , n2899 );
xor ( n5552 , n5312 , n2899 );
xor ( n5553 , n5302 , n2899 );
and ( n5554 , n5487 , n2899 );
and ( n5555 , n5553 , n5554 );
and ( n5556 , n5552 , n5555 );
and ( n5557 , n5551 , n5556 );
and ( n5558 , n5550 , n5557 );
and ( n5559 , n5549 , n5558 );
and ( n5560 , n5548 , n5559 );
and ( n5561 , n5547 , n5560 );
and ( n5562 , n5546 , n5561 );
and ( n5563 , n5545 , n5562 );
and ( n5564 , n5544 , n5563 );
and ( n5565 , n5543 , n5564 );
and ( n5566 , n5542 , n5565 );
and ( n5567 , n5541 , n5566 );
and ( n5568 , n5540 , n5567 );
and ( n5569 , n5539 , n5568 );
and ( n5570 , n5538 , n5569 );
and ( n5571 , n5537 , n5570 );
and ( n5572 , n5536 , n5571 );
xor ( n5573 , n5535 , n5572 );
and ( n5574 , n5573 , n5484 );
or ( n5575 , n5534 , n5574 );
and ( n5576 , n5575 , n5154 );
or ( n5577 , n5532 , n5576 );
not ( n5578 , n5577 );
and ( n5579 , n4083 , n5578 );
and ( n5580 , n2295 , n5290 );
not ( n5581 , n5484 );
and ( n5582 , n5581 , n5472 );
xor ( n5583 , n5536 , n5571 );
and ( n5584 , n5583 , n5484 );
or ( n5585 , n5582 , n5584 );
and ( n5586 , n5585 , n5154 );
or ( n5587 , n5580 , n5586 );
not ( n5588 , n5587 );
and ( n5589 , n4093 , n5588 );
and ( n5590 , n2296 , n5290 );
not ( n5591 , n5484 );
and ( n5592 , n5591 , n5462 );
xor ( n5593 , n5537 , n5570 );
and ( n5594 , n5593 , n5484 );
or ( n5595 , n5592 , n5594 );
and ( n5596 , n5595 , n5154 );
or ( n5597 , n5590 , n5596 );
not ( n5598 , n5597 );
and ( n5599 , n4103 , n5598 );
and ( n5600 , n2297 , n5290 );
not ( n5601 , n5484 );
and ( n5602 , n5601 , n5452 );
xor ( n5603 , n5538 , n5569 );
and ( n5604 , n5603 , n5484 );
or ( n5605 , n5602 , n5604 );
and ( n5606 , n5605 , n5154 );
or ( n5607 , n5600 , n5606 );
not ( n5608 , n5607 );
and ( n5609 , n4113 , n5608 );
and ( n5610 , n2298 , n5290 );
not ( n5611 , n5484 );
and ( n5612 , n5611 , n5442 );
xor ( n5613 , n5539 , n5568 );
and ( n5614 , n5613 , n5484 );
or ( n5615 , n5612 , n5614 );
and ( n5616 , n5615 , n5154 );
or ( n5617 , n5610 , n5616 );
not ( n5618 , n5617 );
and ( n5619 , n4123 , n5618 );
and ( n5620 , n2299 , n5290 );
not ( n5621 , n5484 );
and ( n5622 , n5621 , n5432 );
xor ( n5623 , n5540 , n5567 );
and ( n5624 , n5623 , n5484 );
or ( n5625 , n5622 , n5624 );
and ( n5626 , n5625 , n5154 );
or ( n5627 , n5620 , n5626 );
not ( n5628 , n5627 );
and ( n5629 , n4133 , n5628 );
and ( n5630 , n2300 , n5290 );
not ( n5631 , n5484 );
and ( n5632 , n5631 , n5422 );
xor ( n5633 , n5541 , n5566 );
and ( n5634 , n5633 , n5484 );
or ( n5635 , n5632 , n5634 );
and ( n5636 , n5635 , n5154 );
or ( n5637 , n5630 , n5636 );
not ( n5638 , n5637 );
and ( n5639 , n4143 , n5638 );
and ( n5640 , n2301 , n5290 );
not ( n5641 , n5484 );
and ( n5642 , n5641 , n5412 );
xor ( n5643 , n5542 , n5565 );
and ( n5644 , n5643 , n5484 );
or ( n5645 , n5642 , n5644 );
and ( n5646 , n5645 , n5154 );
or ( n5647 , n5640 , n5646 );
not ( n5648 , n5647 );
and ( n5649 , n4153 , n5648 );
and ( n5650 , n2302 , n5290 );
not ( n5651 , n5484 );
and ( n5652 , n5651 , n5402 );
xor ( n5653 , n5543 , n5564 );
and ( n5654 , n5653 , n5484 );
or ( n5655 , n5652 , n5654 );
and ( n5656 , n5655 , n5154 );
or ( n5657 , n5650 , n5656 );
not ( n5658 , n5657 );
and ( n5659 , n4163 , n5658 );
and ( n5660 , n2303 , n5290 );
not ( n5661 , n5484 );
and ( n5662 , n5661 , n5392 );
xor ( n5663 , n5544 , n5563 );
and ( n5664 , n5663 , n5484 );
or ( n5665 , n5662 , n5664 );
and ( n5666 , n5665 , n5154 );
or ( n5667 , n5660 , n5666 );
not ( n5668 , n5667 );
and ( n5669 , n4173 , n5668 );
and ( n5670 , n2304 , n5290 );
not ( n5671 , n5484 );
and ( n5672 , n5671 , n5382 );
xor ( n5673 , n5545 , n5562 );
and ( n5674 , n5673 , n5484 );
or ( n5675 , n5672 , n5674 );
and ( n5676 , n5675 , n5154 );
or ( n5677 , n5670 , n5676 );
not ( n5678 , n5677 );
and ( n5679 , n4183 , n5678 );
and ( n5680 , n2305 , n5290 );
not ( n5681 , n5484 );
and ( n5682 , n5681 , n5372 );
xor ( n5683 , n5546 , n5561 );
and ( n5684 , n5683 , n5484 );
or ( n5685 , n5682 , n5684 );
and ( n5686 , n5685 , n5154 );
or ( n5687 , n5680 , n5686 );
not ( n5688 , n5687 );
and ( n5689 , n4193 , n5688 );
and ( n5690 , n2306 , n5290 );
not ( n5691 , n5484 );
and ( n5692 , n5691 , n5362 );
xor ( n5693 , n5547 , n5560 );
and ( n5694 , n5693 , n5484 );
or ( n5695 , n5692 , n5694 );
and ( n5696 , n5695 , n5154 );
or ( n5697 , n5690 , n5696 );
not ( n5698 , n5697 );
and ( n5699 , n4203 , n5698 );
and ( n5700 , n2307 , n5290 );
not ( n5701 , n5484 );
and ( n5702 , n5701 , n5352 );
xor ( n5703 , n5548 , n5559 );
and ( n5704 , n5703 , n5484 );
or ( n5705 , n5702 , n5704 );
and ( n5706 , n5705 , n5154 );
or ( n5707 , n5700 , n5706 );
not ( n5708 , n5707 );
and ( n5709 , n4213 , n5708 );
and ( n5710 , n2308 , n5290 );
not ( n5711 , n5484 );
and ( n5712 , n5711 , n5342 );
xor ( n5713 , n5549 , n5558 );
and ( n5714 , n5713 , n5484 );
or ( n5715 , n5712 , n5714 );
and ( n5716 , n5715 , n5154 );
or ( n5717 , n5710 , n5716 );
not ( n5718 , n5717 );
and ( n5719 , n4223 , n5718 );
and ( n5720 , n2309 , n5290 );
not ( n5721 , n5484 );
and ( n5722 , n5721 , n5332 );
xor ( n5723 , n5550 , n5557 );
and ( n5724 , n5723 , n5484 );
or ( n5725 , n5722 , n5724 );
and ( n5726 , n5725 , n5154 );
or ( n5727 , n5720 , n5726 );
not ( n5728 , n5727 );
and ( n5729 , n4233 , n5728 );
and ( n5730 , n2310 , n5290 );
not ( n5731 , n5484 );
and ( n5732 , n5731 , n5322 );
xor ( n5733 , n5551 , n5556 );
and ( n5734 , n5733 , n5484 );
or ( n5735 , n5732 , n5734 );
and ( n5736 , n5735 , n5154 );
or ( n5737 , n5730 , n5736 );
not ( n5738 , n5737 );
and ( n5739 , n4243 , n5738 );
and ( n5740 , n2311 , n5290 );
not ( n5741 , n5484 );
and ( n5742 , n5741 , n5312 );
xor ( n5743 , n5552 , n5555 );
and ( n5744 , n5743 , n5484 );
or ( n5745 , n5742 , n5744 );
and ( n5746 , n5745 , n5154 );
or ( n5747 , n5740 , n5746 );
not ( n5748 , n5747 );
and ( n5749 , n4257 , n5748 );
and ( n5750 , n2312 , n5290 );
not ( n5751 , n5484 );
and ( n5752 , n5751 , n5302 );
xor ( n5753 , n5553 , n5554 );
and ( n5754 , n5753 , n5484 );
or ( n5755 , n5752 , n5754 );
and ( n5756 , n5755 , n5154 );
or ( n5757 , n5750 , n5756 );
not ( n5758 , n5757 );
and ( n5759 , n3785 , n5758 );
not ( n5760 , n5492 );
or ( n5761 , n3795 , n5760 );
and ( n5762 , n5758 , n5761 );
and ( n5763 , n3785 , n5761 );
or ( n5764 , n5759 , n5762 , n5763 );
and ( n5765 , n5748 , n5764 );
and ( n5766 , n4257 , n5764 );
or ( n5767 , n5749 , n5765 , n5766 );
and ( n5768 , n5738 , n5767 );
and ( n5769 , n4243 , n5767 );
or ( n5770 , n5739 , n5768 , n5769 );
and ( n5771 , n5728 , n5770 );
and ( n5772 , n4233 , n5770 );
or ( n5773 , n5729 , n5771 , n5772 );
and ( n5774 , n5718 , n5773 );
and ( n5775 , n4223 , n5773 );
or ( n5776 , n5719 , n5774 , n5775 );
and ( n5777 , n5708 , n5776 );
and ( n5778 , n4213 , n5776 );
or ( n5779 , n5709 , n5777 , n5778 );
and ( n5780 , n5698 , n5779 );
and ( n5781 , n4203 , n5779 );
or ( n5782 , n5699 , n5780 , n5781 );
and ( n5783 , n5688 , n5782 );
and ( n5784 , n4193 , n5782 );
or ( n5785 , n5689 , n5783 , n5784 );
and ( n5786 , n5678 , n5785 );
and ( n5787 , n4183 , n5785 );
or ( n5788 , n5679 , n5786 , n5787 );
and ( n5789 , n5668 , n5788 );
and ( n5790 , n4173 , n5788 );
or ( n5791 , n5669 , n5789 , n5790 );
and ( n5792 , n5658 , n5791 );
and ( n5793 , n4163 , n5791 );
or ( n5794 , n5659 , n5792 , n5793 );
and ( n5795 , n5648 , n5794 );
and ( n5796 , n4153 , n5794 );
or ( n5797 , n5649 , n5795 , n5796 );
and ( n5798 , n5638 , n5797 );
and ( n5799 , n4143 , n5797 );
or ( n5800 , n5639 , n5798 , n5799 );
and ( n5801 , n5628 , n5800 );
and ( n5802 , n4133 , n5800 );
or ( n5803 , n5629 , n5801 , n5802 );
and ( n5804 , n5618 , n5803 );
and ( n5805 , n4123 , n5803 );
or ( n5806 , n5619 , n5804 , n5805 );
and ( n5807 , n5608 , n5806 );
and ( n5808 , n4113 , n5806 );
or ( n5809 , n5609 , n5807 , n5808 );
and ( n5810 , n5598 , n5809 );
and ( n5811 , n4103 , n5809 );
or ( n5812 , n5599 , n5810 , n5811 );
and ( n5813 , n5588 , n5812 );
and ( n5814 , n4093 , n5812 );
or ( n5815 , n5589 , n5813 , n5814 );
and ( n5816 , n5578 , n5815 );
and ( n5817 , n4083 , n5815 );
or ( n5818 , n5579 , n5816 , n5817 );
and ( n5819 , n5530 , n5818 );
and ( n5820 , n4073 , n5818 );
or ( n5821 , n5531 , n5819 , n5820 );
and ( n5822 , n5527 , n5821 );
and ( n5823 , n4063 , n5821 );
or ( n5824 , n5528 , n5822 , n5823 );
and ( n5825 , n5524 , n5824 );
and ( n5826 , n4053 , n5824 );
or ( n5827 , n5525 , n5825 , n5826 );
and ( n5828 , n5521 , n5827 );
and ( n5829 , n4043 , n5827 );
or ( n5830 , n5522 , n5828 , n5829 );
and ( n5831 , n5518 , n5830 );
and ( n5832 , n4033 , n5830 );
or ( n5833 , n5519 , n5831 , n5832 );
and ( n5834 , n5515 , n5833 );
and ( n5835 , n4023 , n5833 );
or ( n5836 , n5516 , n5834 , n5835 );
and ( n5837 , n5512 , n5836 );
and ( n5838 , n4013 , n5836 );
or ( n5839 , n5513 , n5837 , n5838 );
and ( n5840 , n5509 , n5839 );
and ( n5841 , n4003 , n5839 );
or ( n5842 , n5510 , n5840 , n5841 );
and ( n5843 , n5506 , n5842 );
and ( n5844 , n3993 , n5842 );
or ( n5845 , n5507 , n5843 , n5844 );
and ( n5846 , n5503 , n5845 );
and ( n5847 , n3983 , n5845 );
or ( n5848 , n5504 , n5846 , n5847 );
and ( n5849 , n5500 , n5848 );
and ( n5850 , n3819 , n5848 );
or ( n5851 , n5501 , n5849 , n5850 );
xor ( n5852 , n5498 , n5851 );
not ( n5853 , n5852 );
xor ( n5854 , n3785 , n5758 );
xor ( n5855 , n5854 , n5761 );
and ( n5856 , n5853 , n5855 );
not ( n5857 , n5855 );
not ( n5858 , n5493 );
xor ( n5859 , n5857 , n5858 );
and ( n5860 , n5859 , n5852 );
or ( n5861 , n5856 , n5860 );
not ( n5862 , n5861 );
not ( n5863 , n5862 );
or ( n5864 , n5495 , n5863 );
not ( n5865 , n5852 );
xor ( n5866 , n4257 , n5748 );
xor ( n5867 , n5866 , n5764 );
and ( n5868 , n5865 , n5867 );
not ( n5869 , n5867 );
and ( n5870 , n5857 , n5858 );
xor ( n5871 , n5869 , n5870 );
and ( n5872 , n5871 , n5852 );
or ( n5873 , n5868 , n5872 );
not ( n5874 , n5873 );
not ( n5875 , n5874 );
or ( n5876 , n5864 , n5875 );
not ( n5877 , n5852 );
xor ( n5878 , n4243 , n5738 );
xor ( n5879 , n5878 , n5767 );
and ( n5880 , n5877 , n5879 );
not ( n5881 , n5879 );
and ( n5882 , n5869 , n5870 );
xor ( n5883 , n5881 , n5882 );
and ( n5884 , n5883 , n5852 );
or ( n5885 , n5880 , n5884 );
not ( n5886 , n5885 );
not ( n5887 , n5886 );
or ( n5888 , n5876 , n5887 );
not ( n5889 , n5852 );
xor ( n5890 , n4233 , n5728 );
xor ( n5891 , n5890 , n5770 );
and ( n5892 , n5889 , n5891 );
not ( n5893 , n5891 );
and ( n5894 , n5881 , n5882 );
xor ( n5895 , n5893 , n5894 );
and ( n5896 , n5895 , n5852 );
or ( n5897 , n5892 , n5896 );
not ( n5898 , n5897 );
not ( n5899 , n5898 );
or ( n5900 , n5888 , n5899 );
not ( n5901 , n5852 );
xor ( n5902 , n4223 , n5718 );
xor ( n5903 , n5902 , n5773 );
and ( n5904 , n5901 , n5903 );
not ( n5905 , n5903 );
and ( n5906 , n5893 , n5894 );
xor ( n5907 , n5905 , n5906 );
and ( n5908 , n5907 , n5852 );
or ( n5909 , n5904 , n5908 );
not ( n5910 , n5909 );
not ( n5911 , n5910 );
or ( n5912 , n5900 , n5911 );
not ( n5913 , n5852 );
xor ( n5914 , n4213 , n5708 );
xor ( n5915 , n5914 , n5776 );
and ( n5916 , n5913 , n5915 );
not ( n5917 , n5915 );
and ( n5918 , n5905 , n5906 );
xor ( n5919 , n5917 , n5918 );
and ( n5920 , n5919 , n5852 );
or ( n5921 , n5916 , n5920 );
not ( n5922 , n5921 );
not ( n5923 , n5922 );
or ( n5924 , n5912 , n5923 );
not ( n5925 , n5852 );
xor ( n5926 , n4203 , n5698 );
xor ( n5927 , n5926 , n5779 );
and ( n5928 , n5925 , n5927 );
not ( n5929 , n5927 );
and ( n5930 , n5917 , n5918 );
xor ( n5931 , n5929 , n5930 );
and ( n5932 , n5931 , n5852 );
or ( n5933 , n5928 , n5932 );
not ( n5934 , n5933 );
not ( n5935 , n5934 );
or ( n5936 , n5924 , n5935 );
not ( n5937 , n5852 );
xor ( n5938 , n4193 , n5688 );
xor ( n5939 , n5938 , n5782 );
and ( n5940 , n5937 , n5939 );
not ( n5941 , n5939 );
and ( n5942 , n5929 , n5930 );
xor ( n5943 , n5941 , n5942 );
and ( n5944 , n5943 , n5852 );
or ( n5945 , n5940 , n5944 );
not ( n5946 , n5945 );
not ( n5947 , n5946 );
or ( n5948 , n5936 , n5947 );
not ( n5949 , n5852 );
xor ( n5950 , n4183 , n5678 );
xor ( n5951 , n5950 , n5785 );
and ( n5952 , n5949 , n5951 );
not ( n5953 , n5951 );
and ( n5954 , n5941 , n5942 );
xor ( n5955 , n5953 , n5954 );
and ( n5956 , n5955 , n5852 );
or ( n5957 , n5952 , n5956 );
not ( n5958 , n5957 );
not ( n5959 , n5958 );
or ( n5960 , n5948 , n5959 );
not ( n5961 , n5852 );
xor ( n5962 , n4173 , n5668 );
xor ( n5963 , n5962 , n5788 );
and ( n5964 , n5961 , n5963 );
not ( n5965 , n5963 );
and ( n5966 , n5953 , n5954 );
xor ( n5967 , n5965 , n5966 );
and ( n5968 , n5967 , n5852 );
or ( n5969 , n5964 , n5968 );
not ( n5970 , n5969 );
not ( n5971 , n5970 );
or ( n5972 , n5960 , n5971 );
not ( n5973 , n5852 );
xor ( n5974 , n4163 , n5658 );
xor ( n5975 , n5974 , n5791 );
and ( n5976 , n5973 , n5975 );
not ( n5977 , n5975 );
and ( n5978 , n5965 , n5966 );
xor ( n5979 , n5977 , n5978 );
and ( n5980 , n5979 , n5852 );
or ( n5981 , n5976 , n5980 );
not ( n5982 , n5981 );
not ( n5983 , n5982 );
or ( n5984 , n5972 , n5983 );
not ( n5985 , n5852 );
xor ( n5986 , n4153 , n5648 );
xor ( n5987 , n5986 , n5794 );
and ( n5988 , n5985 , n5987 );
not ( n5989 , n5987 );
and ( n5990 , n5977 , n5978 );
xor ( n5991 , n5989 , n5990 );
and ( n5992 , n5991 , n5852 );
or ( n5993 , n5988 , n5992 );
not ( n5994 , n5993 );
not ( n5995 , n5994 );
or ( n5996 , n5984 , n5995 );
not ( n5997 , n5852 );
xor ( n5998 , n4143 , n5638 );
xor ( n5999 , n5998 , n5797 );
and ( n6000 , n5997 , n5999 );
not ( n6001 , n5999 );
and ( n6002 , n5989 , n5990 );
xor ( n6003 , n6001 , n6002 );
and ( n6004 , n6003 , n5852 );
or ( n6005 , n6000 , n6004 );
not ( n6006 , n6005 );
not ( n6007 , n6006 );
or ( n6008 , n5996 , n6007 );
not ( n6009 , n5852 );
xor ( n6010 , n4133 , n5628 );
xor ( n6011 , n6010 , n5800 );
and ( n6012 , n6009 , n6011 );
not ( n6013 , n6011 );
and ( n6014 , n6001 , n6002 );
xor ( n6015 , n6013 , n6014 );
and ( n6016 , n6015 , n5852 );
or ( n6017 , n6012 , n6016 );
not ( n6018 , n6017 );
not ( n6019 , n6018 );
or ( n6020 , n6008 , n6019 );
not ( n6021 , n5852 );
xor ( n6022 , n4123 , n5618 );
xor ( n6023 , n6022 , n5803 );
and ( n6024 , n6021 , n6023 );
not ( n6025 , n6023 );
and ( n6026 , n6013 , n6014 );
xor ( n6027 , n6025 , n6026 );
and ( n6028 , n6027 , n5852 );
or ( n6029 , n6024 , n6028 );
not ( n6030 , n6029 );
not ( n6031 , n6030 );
or ( n6032 , n6020 , n6031 );
not ( n6033 , n5852 );
xor ( n6034 , n4113 , n5608 );
xor ( n6035 , n6034 , n5806 );
and ( n6036 , n6033 , n6035 );
not ( n6037 , n6035 );
and ( n6038 , n6025 , n6026 );
xor ( n6039 , n6037 , n6038 );
and ( n6040 , n6039 , n5852 );
or ( n6041 , n6036 , n6040 );
not ( n6042 , n6041 );
not ( n6043 , n6042 );
or ( n6044 , n6032 , n6043 );
not ( n6045 , n5852 );
xor ( n6046 , n4103 , n5598 );
xor ( n6047 , n6046 , n5809 );
and ( n6048 , n6045 , n6047 );
not ( n6049 , n6047 );
and ( n6050 , n6037 , n6038 );
xor ( n6051 , n6049 , n6050 );
and ( n6052 , n6051 , n5852 );
or ( n6053 , n6048 , n6052 );
not ( n6054 , n6053 );
not ( n6055 , n6054 );
or ( n6056 , n6044 , n6055 );
not ( n6057 , n5852 );
xor ( n6058 , n4093 , n5588 );
xor ( n6059 , n6058 , n5812 );
and ( n6060 , n6057 , n6059 );
not ( n6061 , n6059 );
and ( n6062 , n6049 , n6050 );
xor ( n6063 , n6061 , n6062 );
and ( n6064 , n6063 , n5852 );
or ( n6065 , n6060 , n6064 );
not ( n6066 , n6065 );
not ( n6067 , n6066 );
or ( n6068 , n6056 , n6067 );
not ( n6069 , n5852 );
xor ( n6070 , n4083 , n5578 );
xor ( n6071 , n6070 , n5815 );
and ( n6072 , n6069 , n6071 );
not ( n6073 , n6071 );
and ( n6074 , n6061 , n6062 );
xor ( n6075 , n6073 , n6074 );
and ( n6076 , n6075 , n5852 );
or ( n6077 , n6072 , n6076 );
not ( n6078 , n6077 );
not ( n6079 , n6078 );
or ( n6080 , n6068 , n6079 );
not ( n6081 , n5852 );
xor ( n6082 , n4073 , n5530 );
xor ( n6083 , n6082 , n5818 );
and ( n6084 , n6081 , n6083 );
not ( n6085 , n6083 );
and ( n6086 , n6073 , n6074 );
xor ( n6087 , n6085 , n6086 );
and ( n6088 , n6087 , n5852 );
or ( n6089 , n6084 , n6088 );
not ( n6090 , n6089 );
not ( n6091 , n6090 );
or ( n6092 , n6080 , n6091 );
not ( n6093 , n5852 );
xor ( n6094 , n4063 , n5527 );
xor ( n6095 , n6094 , n5821 );
and ( n6096 , n6093 , n6095 );
not ( n6097 , n6095 );
and ( n6098 , n6085 , n6086 );
xor ( n6099 , n6097 , n6098 );
and ( n6100 , n6099 , n5852 );
or ( n6101 , n6096 , n6100 );
not ( n6102 , n6101 );
not ( n6103 , n6102 );
or ( n6104 , n6092 , n6103 );
not ( n6105 , n5852 );
xor ( n6106 , n4053 , n5524 );
xor ( n6107 , n6106 , n5824 );
and ( n6108 , n6105 , n6107 );
not ( n6109 , n6107 );
and ( n6110 , n6097 , n6098 );
xor ( n6111 , n6109 , n6110 );
and ( n6112 , n6111 , n5852 );
or ( n6113 , n6108 , n6112 );
not ( n6114 , n6113 );
not ( n6115 , n6114 );
or ( n6116 , n6104 , n6115 );
not ( n6117 , n5852 );
xor ( n6118 , n4043 , n5521 );
xor ( n6119 , n6118 , n5827 );
and ( n6120 , n6117 , n6119 );
not ( n6121 , n6119 );
and ( n6122 , n6109 , n6110 );
xor ( n6123 , n6121 , n6122 );
and ( n6124 , n6123 , n5852 );
or ( n6125 , n6120 , n6124 );
not ( n6126 , n6125 );
not ( n6127 , n6126 );
or ( n6128 , n6116 , n6127 );
not ( n6129 , n5852 );
xor ( n6130 , n4033 , n5518 );
xor ( n6131 , n6130 , n5830 );
and ( n6132 , n6129 , n6131 );
not ( n6133 , n6131 );
and ( n6134 , n6121 , n6122 );
xor ( n6135 , n6133 , n6134 );
and ( n6136 , n6135 , n5852 );
or ( n6137 , n6132 , n6136 );
not ( n6138 , n6137 );
not ( n6139 , n6138 );
or ( n6140 , n6128 , n6139 );
not ( n6141 , n5852 );
xor ( n6142 , n4023 , n5515 );
xor ( n6143 , n6142 , n5833 );
and ( n6144 , n6141 , n6143 );
not ( n6145 , n6143 );
and ( n6146 , n6133 , n6134 );
xor ( n6147 , n6145 , n6146 );
and ( n6148 , n6147 , n5852 );
or ( n6149 , n6144 , n6148 );
not ( n6150 , n6149 );
not ( n6151 , n6150 );
or ( n6152 , n6140 , n6151 );
not ( n6153 , n5852 );
xor ( n6154 , n4013 , n5512 );
xor ( n6155 , n6154 , n5836 );
and ( n6156 , n6153 , n6155 );
not ( n6157 , n6155 );
and ( n6158 , n6145 , n6146 );
xor ( n6159 , n6157 , n6158 );
and ( n6160 , n6159 , n5852 );
or ( n6161 , n6156 , n6160 );
not ( n6162 , n6161 );
not ( n6163 , n6162 );
or ( n6164 , n6152 , n6163 );
not ( n6165 , n5852 );
xor ( n6166 , n4003 , n5509 );
xor ( n6167 , n6166 , n5839 );
and ( n6168 , n6165 , n6167 );
not ( n6169 , n6167 );
and ( n6170 , n6157 , n6158 );
xor ( n6171 , n6169 , n6170 );
and ( n6172 , n6171 , n5852 );
or ( n6173 , n6168 , n6172 );
not ( n6174 , n6173 );
not ( n6175 , n6174 );
or ( n6176 , n6164 , n6175 );
not ( n6177 , n5852 );
xor ( n6178 , n3993 , n5506 );
xor ( n6179 , n6178 , n5842 );
and ( n6180 , n6177 , n6179 );
not ( n6181 , n6179 );
and ( n6182 , n6169 , n6170 );
xor ( n6183 , n6181 , n6182 );
and ( n6184 , n6183 , n5852 );
or ( n6185 , n6180 , n6184 );
not ( n6186 , n6185 );
not ( n6187 , n6186 );
or ( n6188 , n6176 , n6187 );
not ( n6189 , n5852 );
xor ( n6190 , n3983 , n5503 );
xor ( n6191 , n6190 , n5845 );
and ( n6192 , n6189 , n6191 );
not ( n6193 , n6191 );
and ( n6194 , n6181 , n6182 );
xor ( n6195 , n6193 , n6194 );
and ( n6196 , n6195 , n5852 );
or ( n6197 , n6192 , n6196 );
not ( n6198 , n6197 );
not ( n6199 , n6198 );
or ( n6200 , n6188 , n6199 );
and ( n6201 , n6200 , n5852 );
not ( n6202 , n6201 );
and ( n6203 , n6202 , n5495 );
xor ( n6204 , n5495 , n5852 );
xor ( n6205 , n6204 , n5852 );
and ( n6206 , n6205 , n6201 );
or ( n6207 , n6203 , n6206 );
and ( n6208 , n6207 , n5188 );
and ( n6209 , n3363 , n5282 );
or ( n6210 , n6208 , n6209 );
not ( n6211 , n3625 );
and ( n6212 , n3627 , n3610 , n3618 , n6211 );
and ( n6213 , n3603 , n3610 , n3618 , n6211 );
or ( n6214 , n6212 , n6213 );
nor ( n6215 , n3627 , n3610 , n3618 , n6211 );
or ( n6216 , n6214 , n6215 );
nor ( n6217 , n3627 , n3611 , n3618 , n6211 );
or ( n6218 , n6216 , n6217 );
and ( n6219 , n6210 , n6218 );
xor ( n6220 , n3795 , n5492 );
not ( n6221 , n6220 );
not ( n6222 , n6221 );
xor ( n6223 , n3770 , n5496 );
and ( n6224 , n3819 , n5499 );
and ( n6225 , n3983 , n5502 );
and ( n6226 , n3993 , n5505 );
and ( n6227 , n4003 , n5508 );
and ( n6228 , n4013 , n5511 );
and ( n6229 , n4023 , n5514 );
and ( n6230 , n4033 , n5517 );
and ( n6231 , n4043 , n5520 );
and ( n6232 , n4053 , n5523 );
and ( n6233 , n4063 , n5526 );
and ( n6234 , n4073 , n5529 );
and ( n6235 , n4083 , n5577 );
and ( n6236 , n4093 , n5587 );
and ( n6237 , n4103 , n5597 );
and ( n6238 , n4113 , n5607 );
and ( n6239 , n4123 , n5617 );
and ( n6240 , n4133 , n5627 );
and ( n6241 , n4143 , n5637 );
and ( n6242 , n4153 , n5647 );
and ( n6243 , n4163 , n5657 );
and ( n6244 , n4173 , n5667 );
and ( n6245 , n4183 , n5677 );
and ( n6246 , n4193 , n5687 );
and ( n6247 , n4203 , n5697 );
and ( n6248 , n4213 , n5707 );
and ( n6249 , n4223 , n5717 );
and ( n6250 , n4233 , n5727 );
and ( n6251 , n4243 , n5737 );
and ( n6252 , n4257 , n5747 );
and ( n6253 , n3785 , n5757 );
and ( n6254 , n3795 , n5492 );
and ( n6255 , n5757 , n6254 );
and ( n6256 , n3785 , n6254 );
or ( n6257 , n6253 , n6255 , n6256 );
and ( n6258 , n5747 , n6257 );
and ( n6259 , n4257 , n6257 );
or ( n6260 , n6252 , n6258 , n6259 );
and ( n6261 , n5737 , n6260 );
and ( n6262 , n4243 , n6260 );
or ( n6263 , n6251 , n6261 , n6262 );
and ( n6264 , n5727 , n6263 );
and ( n6265 , n4233 , n6263 );
or ( n6266 , n6250 , n6264 , n6265 );
and ( n6267 , n5717 , n6266 );
and ( n6268 , n4223 , n6266 );
or ( n6269 , n6249 , n6267 , n6268 );
and ( n6270 , n5707 , n6269 );
and ( n6271 , n4213 , n6269 );
or ( n6272 , n6248 , n6270 , n6271 );
and ( n6273 , n5697 , n6272 );
and ( n6274 , n4203 , n6272 );
or ( n6275 , n6247 , n6273 , n6274 );
and ( n6276 , n5687 , n6275 );
and ( n6277 , n4193 , n6275 );
or ( n6278 , n6246 , n6276 , n6277 );
and ( n6279 , n5677 , n6278 );
and ( n6280 , n4183 , n6278 );
or ( n6281 , n6245 , n6279 , n6280 );
and ( n6282 , n5667 , n6281 );
and ( n6283 , n4173 , n6281 );
or ( n6284 , n6244 , n6282 , n6283 );
and ( n6285 , n5657 , n6284 );
and ( n6286 , n4163 , n6284 );
or ( n6287 , n6243 , n6285 , n6286 );
and ( n6288 , n5647 , n6287 );
and ( n6289 , n4153 , n6287 );
or ( n6290 , n6242 , n6288 , n6289 );
and ( n6291 , n5637 , n6290 );
and ( n6292 , n4143 , n6290 );
or ( n6293 , n6241 , n6291 , n6292 );
and ( n6294 , n5627 , n6293 );
and ( n6295 , n4133 , n6293 );
or ( n6296 , n6240 , n6294 , n6295 );
and ( n6297 , n5617 , n6296 );
and ( n6298 , n4123 , n6296 );
or ( n6299 , n6239 , n6297 , n6298 );
and ( n6300 , n5607 , n6299 );
and ( n6301 , n4113 , n6299 );
or ( n6302 , n6238 , n6300 , n6301 );
and ( n6303 , n5597 , n6302 );
and ( n6304 , n4103 , n6302 );
or ( n6305 , n6237 , n6303 , n6304 );
and ( n6306 , n5587 , n6305 );
and ( n6307 , n4093 , n6305 );
or ( n6308 , n6236 , n6306 , n6307 );
and ( n6309 , n5577 , n6308 );
and ( n6310 , n4083 , n6308 );
or ( n6311 , n6235 , n6309 , n6310 );
and ( n6312 , n5529 , n6311 );
and ( n6313 , n4073 , n6311 );
or ( n6314 , n6234 , n6312 , n6313 );
and ( n6315 , n5526 , n6314 );
and ( n6316 , n4063 , n6314 );
or ( n6317 , n6233 , n6315 , n6316 );
and ( n6318 , n5523 , n6317 );
and ( n6319 , n4053 , n6317 );
or ( n6320 , n6232 , n6318 , n6319 );
and ( n6321 , n5520 , n6320 );
and ( n6322 , n4043 , n6320 );
or ( n6323 , n6231 , n6321 , n6322 );
and ( n6324 , n5517 , n6323 );
and ( n6325 , n4033 , n6323 );
or ( n6326 , n6230 , n6324 , n6325 );
and ( n6327 , n5514 , n6326 );
and ( n6328 , n4023 , n6326 );
or ( n6329 , n6229 , n6327 , n6328 );
and ( n6330 , n5511 , n6329 );
and ( n6331 , n4013 , n6329 );
or ( n6332 , n6228 , n6330 , n6331 );
and ( n6333 , n5508 , n6332 );
and ( n6334 , n4003 , n6332 );
or ( n6335 , n6227 , n6333 , n6334 );
and ( n6336 , n5505 , n6335 );
and ( n6337 , n3993 , n6335 );
or ( n6338 , n6226 , n6336 , n6337 );
and ( n6339 , n5502 , n6338 );
and ( n6340 , n3983 , n6338 );
or ( n6341 , n6225 , n6339 , n6340 );
and ( n6342 , n5499 , n6341 );
and ( n6343 , n3819 , n6341 );
or ( n6344 , n6224 , n6342 , n6343 );
xor ( n6345 , n6223 , n6344 );
not ( n6346 , n6345 );
xor ( n6347 , n3785 , n5757 );
xor ( n6348 , n6347 , n6254 );
and ( n6349 , n6346 , n6348 );
not ( n6350 , n6348 );
not ( n6351 , n6220 );
xor ( n6352 , n6350 , n6351 );
and ( n6353 , n6352 , n6345 );
or ( n6354 , n6349 , n6353 );
not ( n6355 , n6354 );
not ( n6356 , n6355 );
or ( n6357 , n6222 , n6356 );
not ( n6358 , n6345 );
xor ( n6359 , n4257 , n5747 );
xor ( n6360 , n6359 , n6257 );
and ( n6361 , n6358 , n6360 );
not ( n6362 , n6360 );
and ( n6363 , n6350 , n6351 );
xor ( n6364 , n6362 , n6363 );
and ( n6365 , n6364 , n6345 );
or ( n6366 , n6361 , n6365 );
not ( n6367 , n6366 );
not ( n6368 , n6367 );
or ( n6369 , n6357 , n6368 );
not ( n6370 , n6345 );
xor ( n6371 , n4243 , n5737 );
xor ( n6372 , n6371 , n6260 );
and ( n6373 , n6370 , n6372 );
not ( n6374 , n6372 );
and ( n6375 , n6362 , n6363 );
xor ( n6376 , n6374 , n6375 );
and ( n6377 , n6376 , n6345 );
or ( n6378 , n6373 , n6377 );
not ( n6379 , n6378 );
not ( n6380 , n6379 );
or ( n6381 , n6369 , n6380 );
not ( n6382 , n6345 );
xor ( n6383 , n4233 , n5727 );
xor ( n6384 , n6383 , n6263 );
and ( n6385 , n6382 , n6384 );
not ( n6386 , n6384 );
and ( n6387 , n6374 , n6375 );
xor ( n6388 , n6386 , n6387 );
and ( n6389 , n6388 , n6345 );
or ( n6390 , n6385 , n6389 );
not ( n6391 , n6390 );
not ( n6392 , n6391 );
or ( n6393 , n6381 , n6392 );
not ( n6394 , n6345 );
xor ( n6395 , n4223 , n5717 );
xor ( n6396 , n6395 , n6266 );
and ( n6397 , n6394 , n6396 );
not ( n6398 , n6396 );
and ( n6399 , n6386 , n6387 );
xor ( n6400 , n6398 , n6399 );
and ( n6401 , n6400 , n6345 );
or ( n6402 , n6397 , n6401 );
not ( n6403 , n6402 );
not ( n6404 , n6403 );
or ( n6405 , n6393 , n6404 );
not ( n6406 , n6345 );
xor ( n6407 , n4213 , n5707 );
xor ( n6408 , n6407 , n6269 );
and ( n6409 , n6406 , n6408 );
not ( n6410 , n6408 );
and ( n6411 , n6398 , n6399 );
xor ( n6412 , n6410 , n6411 );
and ( n6413 , n6412 , n6345 );
or ( n6414 , n6409 , n6413 );
not ( n6415 , n6414 );
not ( n6416 , n6415 );
or ( n6417 , n6405 , n6416 );
not ( n6418 , n6345 );
xor ( n6419 , n4203 , n5697 );
xor ( n6420 , n6419 , n6272 );
and ( n6421 , n6418 , n6420 );
not ( n6422 , n6420 );
and ( n6423 , n6410 , n6411 );
xor ( n6424 , n6422 , n6423 );
and ( n6425 , n6424 , n6345 );
or ( n6426 , n6421 , n6425 );
not ( n6427 , n6426 );
not ( n6428 , n6427 );
or ( n6429 , n6417 , n6428 );
not ( n6430 , n6345 );
xor ( n6431 , n4193 , n5687 );
xor ( n6432 , n6431 , n6275 );
and ( n6433 , n6430 , n6432 );
not ( n6434 , n6432 );
and ( n6435 , n6422 , n6423 );
xor ( n6436 , n6434 , n6435 );
and ( n6437 , n6436 , n6345 );
or ( n6438 , n6433 , n6437 );
not ( n6439 , n6438 );
not ( n6440 , n6439 );
or ( n6441 , n6429 , n6440 );
not ( n6442 , n6345 );
xor ( n6443 , n4183 , n5677 );
xor ( n6444 , n6443 , n6278 );
and ( n6445 , n6442 , n6444 );
not ( n6446 , n6444 );
and ( n6447 , n6434 , n6435 );
xor ( n6448 , n6446 , n6447 );
and ( n6449 , n6448 , n6345 );
or ( n6450 , n6445 , n6449 );
not ( n6451 , n6450 );
not ( n6452 , n6451 );
or ( n6453 , n6441 , n6452 );
not ( n6454 , n6345 );
xor ( n6455 , n4173 , n5667 );
xor ( n6456 , n6455 , n6281 );
and ( n6457 , n6454 , n6456 );
not ( n6458 , n6456 );
and ( n6459 , n6446 , n6447 );
xor ( n6460 , n6458 , n6459 );
and ( n6461 , n6460 , n6345 );
or ( n6462 , n6457 , n6461 );
not ( n6463 , n6462 );
not ( n6464 , n6463 );
or ( n6465 , n6453 , n6464 );
not ( n6466 , n6345 );
xor ( n6467 , n4163 , n5657 );
xor ( n6468 , n6467 , n6284 );
and ( n6469 , n6466 , n6468 );
not ( n6470 , n6468 );
and ( n6471 , n6458 , n6459 );
xor ( n6472 , n6470 , n6471 );
and ( n6473 , n6472 , n6345 );
or ( n6474 , n6469 , n6473 );
not ( n6475 , n6474 );
not ( n6476 , n6475 );
or ( n6477 , n6465 , n6476 );
not ( n6478 , n6345 );
xor ( n6479 , n4153 , n5647 );
xor ( n6480 , n6479 , n6287 );
and ( n6481 , n6478 , n6480 );
not ( n6482 , n6480 );
and ( n6483 , n6470 , n6471 );
xor ( n6484 , n6482 , n6483 );
and ( n6485 , n6484 , n6345 );
or ( n6486 , n6481 , n6485 );
not ( n6487 , n6486 );
not ( n6488 , n6487 );
or ( n6489 , n6477 , n6488 );
not ( n6490 , n6345 );
xor ( n6491 , n4143 , n5637 );
xor ( n6492 , n6491 , n6290 );
and ( n6493 , n6490 , n6492 );
not ( n6494 , n6492 );
and ( n6495 , n6482 , n6483 );
xor ( n6496 , n6494 , n6495 );
and ( n6497 , n6496 , n6345 );
or ( n6498 , n6493 , n6497 );
not ( n6499 , n6498 );
not ( n6500 , n6499 );
or ( n6501 , n6489 , n6500 );
not ( n6502 , n6345 );
xor ( n6503 , n4133 , n5627 );
xor ( n6504 , n6503 , n6293 );
and ( n6505 , n6502 , n6504 );
not ( n6506 , n6504 );
and ( n6507 , n6494 , n6495 );
xor ( n6508 , n6506 , n6507 );
and ( n6509 , n6508 , n6345 );
or ( n6510 , n6505 , n6509 );
not ( n6511 , n6510 );
not ( n6512 , n6511 );
or ( n6513 , n6501 , n6512 );
not ( n6514 , n6345 );
xor ( n6515 , n4123 , n5617 );
xor ( n6516 , n6515 , n6296 );
and ( n6517 , n6514 , n6516 );
not ( n6518 , n6516 );
and ( n6519 , n6506 , n6507 );
xor ( n6520 , n6518 , n6519 );
and ( n6521 , n6520 , n6345 );
or ( n6522 , n6517 , n6521 );
not ( n6523 , n6522 );
not ( n6524 , n6523 );
or ( n6525 , n6513 , n6524 );
not ( n6526 , n6345 );
xor ( n6527 , n4113 , n5607 );
xor ( n6528 , n6527 , n6299 );
and ( n6529 , n6526 , n6528 );
not ( n6530 , n6528 );
and ( n6531 , n6518 , n6519 );
xor ( n6532 , n6530 , n6531 );
and ( n6533 , n6532 , n6345 );
or ( n6534 , n6529 , n6533 );
not ( n6535 , n6534 );
not ( n6536 , n6535 );
or ( n6537 , n6525 , n6536 );
not ( n6538 , n6345 );
xor ( n6539 , n4103 , n5597 );
xor ( n6540 , n6539 , n6302 );
and ( n6541 , n6538 , n6540 );
not ( n6542 , n6540 );
and ( n6543 , n6530 , n6531 );
xor ( n6544 , n6542 , n6543 );
and ( n6545 , n6544 , n6345 );
or ( n6546 , n6541 , n6545 );
not ( n6547 , n6546 );
not ( n6548 , n6547 );
or ( n6549 , n6537 , n6548 );
not ( n6550 , n6345 );
xor ( n6551 , n4093 , n5587 );
xor ( n6552 , n6551 , n6305 );
and ( n6553 , n6550 , n6552 );
not ( n6554 , n6552 );
and ( n6555 , n6542 , n6543 );
xor ( n6556 , n6554 , n6555 );
and ( n6557 , n6556 , n6345 );
or ( n6558 , n6553 , n6557 );
not ( n6559 , n6558 );
not ( n6560 , n6559 );
or ( n6561 , n6549 , n6560 );
not ( n6562 , n6345 );
xor ( n6563 , n4083 , n5577 );
xor ( n6564 , n6563 , n6308 );
and ( n6565 , n6562 , n6564 );
not ( n6566 , n6564 );
and ( n6567 , n6554 , n6555 );
xor ( n6568 , n6566 , n6567 );
and ( n6569 , n6568 , n6345 );
or ( n6570 , n6565 , n6569 );
not ( n6571 , n6570 );
not ( n6572 , n6571 );
or ( n6573 , n6561 , n6572 );
not ( n6574 , n6345 );
xor ( n6575 , n4073 , n5529 );
xor ( n6576 , n6575 , n6311 );
and ( n6577 , n6574 , n6576 );
not ( n6578 , n6576 );
and ( n6579 , n6566 , n6567 );
xor ( n6580 , n6578 , n6579 );
and ( n6581 , n6580 , n6345 );
or ( n6582 , n6577 , n6581 );
not ( n6583 , n6582 );
not ( n6584 , n6583 );
or ( n6585 , n6573 , n6584 );
not ( n6586 , n6345 );
xor ( n6587 , n4063 , n5526 );
xor ( n6588 , n6587 , n6314 );
and ( n6589 , n6586 , n6588 );
not ( n6590 , n6588 );
and ( n6591 , n6578 , n6579 );
xor ( n6592 , n6590 , n6591 );
and ( n6593 , n6592 , n6345 );
or ( n6594 , n6589 , n6593 );
not ( n6595 , n6594 );
not ( n6596 , n6595 );
or ( n6597 , n6585 , n6596 );
not ( n6598 , n6345 );
xor ( n6599 , n4053 , n5523 );
xor ( n6600 , n6599 , n6317 );
and ( n6601 , n6598 , n6600 );
not ( n6602 , n6600 );
and ( n6603 , n6590 , n6591 );
xor ( n6604 , n6602 , n6603 );
and ( n6605 , n6604 , n6345 );
or ( n6606 , n6601 , n6605 );
not ( n6607 , n6606 );
not ( n6608 , n6607 );
or ( n6609 , n6597 , n6608 );
not ( n6610 , n6345 );
xor ( n6611 , n4043 , n5520 );
xor ( n6612 , n6611 , n6320 );
and ( n6613 , n6610 , n6612 );
not ( n6614 , n6612 );
and ( n6615 , n6602 , n6603 );
xor ( n6616 , n6614 , n6615 );
and ( n6617 , n6616 , n6345 );
or ( n6618 , n6613 , n6617 );
not ( n6619 , n6618 );
not ( n6620 , n6619 );
or ( n6621 , n6609 , n6620 );
not ( n6622 , n6345 );
xor ( n6623 , n4033 , n5517 );
xor ( n6624 , n6623 , n6323 );
and ( n6625 , n6622 , n6624 );
not ( n6626 , n6624 );
and ( n6627 , n6614 , n6615 );
xor ( n6628 , n6626 , n6627 );
and ( n6629 , n6628 , n6345 );
or ( n6630 , n6625 , n6629 );
not ( n6631 , n6630 );
not ( n6632 , n6631 );
or ( n6633 , n6621 , n6632 );
not ( n6634 , n6345 );
xor ( n6635 , n4023 , n5514 );
xor ( n6636 , n6635 , n6326 );
and ( n6637 , n6634 , n6636 );
not ( n6638 , n6636 );
and ( n6639 , n6626 , n6627 );
xor ( n6640 , n6638 , n6639 );
and ( n6641 , n6640 , n6345 );
or ( n6642 , n6637 , n6641 );
not ( n6643 , n6642 );
not ( n6644 , n6643 );
or ( n6645 , n6633 , n6644 );
not ( n6646 , n6345 );
xor ( n6647 , n4013 , n5511 );
xor ( n6648 , n6647 , n6329 );
and ( n6649 , n6646 , n6648 );
not ( n6650 , n6648 );
and ( n6651 , n6638 , n6639 );
xor ( n6652 , n6650 , n6651 );
and ( n6653 , n6652 , n6345 );
or ( n6654 , n6649 , n6653 );
not ( n6655 , n6654 );
not ( n6656 , n6655 );
or ( n6657 , n6645 , n6656 );
not ( n6658 , n6345 );
xor ( n6659 , n4003 , n5508 );
xor ( n6660 , n6659 , n6332 );
and ( n6661 , n6658 , n6660 );
not ( n6662 , n6660 );
and ( n6663 , n6650 , n6651 );
xor ( n6664 , n6662 , n6663 );
and ( n6665 , n6664 , n6345 );
or ( n6666 , n6661 , n6665 );
not ( n6667 , n6666 );
not ( n6668 , n6667 );
or ( n6669 , n6657 , n6668 );
not ( n6670 , n6345 );
xor ( n6671 , n3993 , n5505 );
xor ( n6672 , n6671 , n6335 );
and ( n6673 , n6670 , n6672 );
not ( n6674 , n6672 );
and ( n6675 , n6662 , n6663 );
xor ( n6676 , n6674 , n6675 );
and ( n6677 , n6676 , n6345 );
or ( n6678 , n6673 , n6677 );
not ( n6679 , n6678 );
not ( n6680 , n6679 );
or ( n6681 , n6669 , n6680 );
not ( n6682 , n6345 );
xor ( n6683 , n3983 , n5502 );
xor ( n6684 , n6683 , n6338 );
and ( n6685 , n6682 , n6684 );
not ( n6686 , n6684 );
and ( n6687 , n6674 , n6675 );
xor ( n6688 , n6686 , n6687 );
and ( n6689 , n6688 , n6345 );
or ( n6690 , n6685 , n6689 );
not ( n6691 , n6690 );
not ( n6692 , n6691 );
or ( n6693 , n6681 , n6692 );
and ( n6694 , n6693 , n6345 );
not ( n6695 , n6694 );
and ( n6696 , n6695 , n6222 );
xor ( n6697 , n6222 , n6345 );
xor ( n6698 , n6697 , n6345 );
and ( n6699 , n6698 , n6694 );
or ( n6700 , n6696 , n6699 );
and ( n6701 , n6700 , n5188 );
and ( n6702 , n3363 , n5282 );
or ( n6703 , n6701 , n6702 );
and ( n6704 , n3627 , n3611 , n3618 , n6211 );
and ( n6705 , n3603 , n3611 , n3618 , n6211 );
or ( n6706 , n6704 , n6705 );
nor ( n6707 , n3603 , n3610 , n3618 , n6211 );
or ( n6708 , n6706 , n6707 );
nor ( n6709 , n3603 , n3611 , n3618 , n6211 );
or ( n6710 , n6708 , n6709 );
and ( n6711 , n6703 , n6710 );
and ( n6712 , n5492 , n5188 );
and ( n6713 , n3363 , n5282 );
or ( n6714 , n6712 , n6713 );
nor ( n6715 , n3603 , n3611 , n3618 , n3625 );
nor ( n6716 , n3627 , n3611 , n3618 , n3625 );
or ( n6717 , n6715 , n6716 );
and ( n6718 , n6714 , n6717 );
nor ( n6719 , n3627 , n3610 , n3618 , n3625 );
and ( n6720 , n5492 , n6719 );
and ( n6721 , n5492 , n5188 );
and ( n6722 , n3363 , n5282 );
or ( n6723 , n6721 , n6722 );
nor ( n6724 , n3603 , n3610 , n3618 , n3625 );
and ( n6725 , n6723 , n6724 );
or ( n6726 , n3632 , n5286 , n6219 , n6711 , n6718 , n6720 , n6725 );
and ( n6727 , n3360 , n6726 );
and ( n6728 , n3363 , n3260 );
or ( n6729 , n6727 , n6728 );
and ( n6730 , n6729 , n2422 );
and ( n6731 , n3356 , n2428 );
or ( n6732 , n6730 , n6731 );
buf ( n6733 , n6732 );
buf ( n6734 , n2424 );
buf ( n6735 , n2281 );
buf ( n6736 , n2280 );
not ( n6737 , n3260 );
and ( n6738 , n3776 , n3631 );
not ( n6739 , n3795 );
not ( n6740 , n6739 );
not ( n6741 , n3770 );
and ( n6742 , n6741 , n3785 );
not ( n6743 , n3785 );
not ( n6744 , n3795 );
xor ( n6745 , n6743 , n6744 );
and ( n6746 , n6745 , n3770 );
or ( n6747 , n6742 , n6746 );
not ( n6748 , n6747 );
not ( n6749 , n6748 );
or ( n6750 , n6740 , n6749 );
not ( n6751 , n3770 );
and ( n6752 , n6751 , n4257 );
not ( n6753 , n4257 );
and ( n6754 , n6743 , n6744 );
xor ( n6755 , n6753 , n6754 );
and ( n6756 , n6755 , n3770 );
or ( n6757 , n6752 , n6756 );
not ( n6758 , n6757 );
not ( n6759 , n6758 );
or ( n6760 , n6750 , n6759 );
not ( n6761 , n3770 );
and ( n6762 , n6761 , n4243 );
not ( n6763 , n4243 );
and ( n6764 , n6753 , n6754 );
xor ( n6765 , n6763 , n6764 );
and ( n6766 , n6765 , n3770 );
or ( n6767 , n6762 , n6766 );
not ( n6768 , n6767 );
not ( n6769 , n6768 );
or ( n6770 , n6760 , n6769 );
not ( n6771 , n3770 );
and ( n6772 , n6771 , n4233 );
not ( n6773 , n4233 );
and ( n6774 , n6763 , n6764 );
xor ( n6775 , n6773 , n6774 );
and ( n6776 , n6775 , n3770 );
or ( n6777 , n6772 , n6776 );
not ( n6778 , n6777 );
not ( n6779 , n6778 );
or ( n6780 , n6770 , n6779 );
not ( n6781 , n3770 );
and ( n6782 , n6781 , n4223 );
not ( n6783 , n4223 );
and ( n6784 , n6773 , n6774 );
xor ( n6785 , n6783 , n6784 );
and ( n6786 , n6785 , n3770 );
or ( n6787 , n6782 , n6786 );
not ( n6788 , n6787 );
not ( n6789 , n6788 );
or ( n6790 , n6780 , n6789 );
not ( n6791 , n3770 );
and ( n6792 , n6791 , n4213 );
not ( n6793 , n4213 );
and ( n6794 , n6783 , n6784 );
xor ( n6795 , n6793 , n6794 );
and ( n6796 , n6795 , n3770 );
or ( n6797 , n6792 , n6796 );
not ( n6798 , n6797 );
not ( n6799 , n6798 );
or ( n6800 , n6790 , n6799 );
not ( n6801 , n3770 );
and ( n6802 , n6801 , n4203 );
not ( n6803 , n4203 );
and ( n6804 , n6793 , n6794 );
xor ( n6805 , n6803 , n6804 );
and ( n6806 , n6805 , n3770 );
or ( n6807 , n6802 , n6806 );
not ( n6808 , n6807 );
not ( n6809 , n6808 );
or ( n6810 , n6800 , n6809 );
not ( n6811 , n3770 );
and ( n6812 , n6811 , n4193 );
not ( n6813 , n4193 );
and ( n6814 , n6803 , n6804 );
xor ( n6815 , n6813 , n6814 );
and ( n6816 , n6815 , n3770 );
or ( n6817 , n6812 , n6816 );
not ( n6818 , n6817 );
not ( n6819 , n6818 );
or ( n6820 , n6810 , n6819 );
not ( n6821 , n3770 );
and ( n6822 , n6821 , n4183 );
not ( n6823 , n4183 );
and ( n6824 , n6813 , n6814 );
xor ( n6825 , n6823 , n6824 );
and ( n6826 , n6825 , n3770 );
or ( n6827 , n6822 , n6826 );
not ( n6828 , n6827 );
not ( n6829 , n6828 );
or ( n6830 , n6820 , n6829 );
not ( n6831 , n3770 );
and ( n6832 , n6831 , n4173 );
not ( n6833 , n4173 );
and ( n6834 , n6823 , n6824 );
xor ( n6835 , n6833 , n6834 );
and ( n6836 , n6835 , n3770 );
or ( n6837 , n6832 , n6836 );
not ( n6838 , n6837 );
not ( n6839 , n6838 );
or ( n6840 , n6830 , n6839 );
not ( n6841 , n3770 );
and ( n6842 , n6841 , n4163 );
not ( n6843 , n4163 );
and ( n6844 , n6833 , n6834 );
xor ( n6845 , n6843 , n6844 );
and ( n6846 , n6845 , n3770 );
or ( n6847 , n6842 , n6846 );
not ( n6848 , n6847 );
not ( n6849 , n6848 );
or ( n6850 , n6840 , n6849 );
not ( n6851 , n3770 );
and ( n6852 , n6851 , n4153 );
not ( n6853 , n4153 );
and ( n6854 , n6843 , n6844 );
xor ( n6855 , n6853 , n6854 );
and ( n6856 , n6855 , n3770 );
or ( n6857 , n6852 , n6856 );
not ( n6858 , n6857 );
not ( n6859 , n6858 );
or ( n6860 , n6850 , n6859 );
not ( n6861 , n3770 );
and ( n6862 , n6861 , n4143 );
not ( n6863 , n4143 );
and ( n6864 , n6853 , n6854 );
xor ( n6865 , n6863 , n6864 );
and ( n6866 , n6865 , n3770 );
or ( n6867 , n6862 , n6866 );
not ( n6868 , n6867 );
not ( n6869 , n6868 );
or ( n6870 , n6860 , n6869 );
not ( n6871 , n3770 );
and ( n6872 , n6871 , n4133 );
not ( n6873 , n4133 );
and ( n6874 , n6863 , n6864 );
xor ( n6875 , n6873 , n6874 );
and ( n6876 , n6875 , n3770 );
or ( n6877 , n6872 , n6876 );
not ( n6878 , n6877 );
not ( n6879 , n6878 );
or ( n6880 , n6870 , n6879 );
not ( n6881 , n3770 );
and ( n6882 , n6881 , n4123 );
not ( n6883 , n4123 );
and ( n6884 , n6873 , n6874 );
xor ( n6885 , n6883 , n6884 );
and ( n6886 , n6885 , n3770 );
or ( n6887 , n6882 , n6886 );
not ( n6888 , n6887 );
not ( n6889 , n6888 );
or ( n6890 , n6880 , n6889 );
not ( n6891 , n3770 );
and ( n6892 , n6891 , n4113 );
not ( n6893 , n4113 );
and ( n6894 , n6883 , n6884 );
xor ( n6895 , n6893 , n6894 );
and ( n6896 , n6895 , n3770 );
or ( n6897 , n6892 , n6896 );
not ( n6898 , n6897 );
not ( n6899 , n6898 );
or ( n6900 , n6890 , n6899 );
not ( n6901 , n3770 );
and ( n6902 , n6901 , n4103 );
not ( n6903 , n4103 );
and ( n6904 , n6893 , n6894 );
xor ( n6905 , n6903 , n6904 );
and ( n6906 , n6905 , n3770 );
or ( n6907 , n6902 , n6906 );
not ( n6908 , n6907 );
not ( n6909 , n6908 );
or ( n6910 , n6900 , n6909 );
not ( n6911 , n3770 );
and ( n6912 , n6911 , n4093 );
not ( n6913 , n4093 );
and ( n6914 , n6903 , n6904 );
xor ( n6915 , n6913 , n6914 );
and ( n6916 , n6915 , n3770 );
or ( n6917 , n6912 , n6916 );
not ( n6918 , n6917 );
not ( n6919 , n6918 );
or ( n6920 , n6910 , n6919 );
not ( n6921 , n3770 );
and ( n6922 , n6921 , n4083 );
not ( n6923 , n4083 );
and ( n6924 , n6913 , n6914 );
xor ( n6925 , n6923 , n6924 );
and ( n6926 , n6925 , n3770 );
or ( n6927 , n6922 , n6926 );
not ( n6928 , n6927 );
not ( n6929 , n6928 );
or ( n6930 , n6920 , n6929 );
not ( n6931 , n3770 );
and ( n6932 , n6931 , n4073 );
not ( n6933 , n4073 );
and ( n6934 , n6923 , n6924 );
xor ( n6935 , n6933 , n6934 );
and ( n6936 , n6935 , n3770 );
or ( n6937 , n6932 , n6936 );
not ( n6938 , n6937 );
not ( n6939 , n6938 );
or ( n6940 , n6930 , n6939 );
not ( n6941 , n3770 );
and ( n6942 , n6941 , n4063 );
not ( n6943 , n4063 );
and ( n6944 , n6933 , n6934 );
xor ( n6945 , n6943 , n6944 );
and ( n6946 , n6945 , n3770 );
or ( n6947 , n6942 , n6946 );
not ( n6948 , n6947 );
not ( n6949 , n6948 );
or ( n6950 , n6940 , n6949 );
not ( n6951 , n3770 );
and ( n6952 , n6951 , n4053 );
not ( n6953 , n4053 );
and ( n6954 , n6943 , n6944 );
xor ( n6955 , n6953 , n6954 );
and ( n6956 , n6955 , n3770 );
or ( n6957 , n6952 , n6956 );
not ( n6958 , n6957 );
not ( n6959 , n6958 );
or ( n6960 , n6950 , n6959 );
not ( n6961 , n3770 );
and ( n6962 , n6961 , n4043 );
not ( n6963 , n4043 );
and ( n6964 , n6953 , n6954 );
xor ( n6965 , n6963 , n6964 );
and ( n6966 , n6965 , n3770 );
or ( n6967 , n6962 , n6966 );
not ( n6968 , n6967 );
not ( n6969 , n6968 );
or ( n6970 , n6960 , n6969 );
not ( n6971 , n3770 );
and ( n6972 , n6971 , n4033 );
not ( n6973 , n4033 );
and ( n6974 , n6963 , n6964 );
xor ( n6975 , n6973 , n6974 );
and ( n6976 , n6975 , n3770 );
or ( n6977 , n6972 , n6976 );
not ( n6978 , n6977 );
not ( n6979 , n6978 );
or ( n6980 , n6970 , n6979 );
not ( n6981 , n3770 );
and ( n6982 , n6981 , n4023 );
not ( n6983 , n4023 );
and ( n6984 , n6973 , n6974 );
xor ( n6985 , n6983 , n6984 );
and ( n6986 , n6985 , n3770 );
or ( n6987 , n6982 , n6986 );
not ( n6988 , n6987 );
not ( n6989 , n6988 );
or ( n6990 , n6980 , n6989 );
not ( n6991 , n3770 );
and ( n6992 , n6991 , n4013 );
not ( n6993 , n4013 );
and ( n6994 , n6983 , n6984 );
xor ( n6995 , n6993 , n6994 );
and ( n6996 , n6995 , n3770 );
or ( n6997 , n6992 , n6996 );
not ( n6998 , n6997 );
not ( n6999 , n6998 );
or ( n7000 , n6990 , n6999 );
not ( n7001 , n3770 );
and ( n7002 , n7001 , n4003 );
not ( n7003 , n4003 );
and ( n7004 , n6993 , n6994 );
xor ( n7005 , n7003 , n7004 );
and ( n7006 , n7005 , n3770 );
or ( n7007 , n7002 , n7006 );
not ( n7008 , n7007 );
not ( n7009 , n7008 );
or ( n7010 , n7000 , n7009 );
not ( n7011 , n3770 );
and ( n7012 , n7011 , n3993 );
not ( n7013 , n3993 );
and ( n7014 , n7003 , n7004 );
xor ( n7015 , n7013 , n7014 );
and ( n7016 , n7015 , n3770 );
or ( n7017 , n7012 , n7016 );
not ( n7018 , n7017 );
not ( n7019 , n7018 );
or ( n7020 , n7010 , n7019 );
and ( n7021 , n7020 , n3770 );
not ( n7022 , n7021 );
and ( n7023 , n7022 , n6740 );
xor ( n7024 , n6740 , n3770 );
xor ( n7025 , n7024 , n3770 );
and ( n7026 , n7025 , n7021 );
or ( n7027 , n7023 , n7026 );
and ( n7028 , n7027 , n5289 );
and ( n7029 , n7027 , n5287 );
not ( n7030 , n3290 );
and ( n7031 , n7030 , n4584 );
not ( n7032 , n4999 );
and ( n7033 , n7032 , n4592 );
xor ( n7034 , n4592 , n4578 );
and ( n7035 , n5002 , n4578 );
xor ( n7036 , n7034 , n7035 );
and ( n7037 , n7036 , n4999 );
or ( n7038 , n7033 , n7037 );
and ( n7039 , n7038 , n3290 );
or ( n7040 , n7031 , n7039 );
and ( n7041 , n7040 , n5152 );
and ( n7042 , n4584 , n5154 );
or ( n7043 , n7028 , n7029 , n7041 , n7042 );
and ( n7044 , n7043 , n5188 );
and ( n7045 , n3776 , n5282 );
or ( n7046 , n7044 , n7045 );
and ( n7047 , n7046 , n5285 );
not ( n7048 , n6201 );
and ( n7049 , n7048 , n5863 );
xor ( n7050 , n5863 , n5852 );
and ( n7051 , n6204 , n5852 );
xor ( n7052 , n7050 , n7051 );
and ( n7053 , n7052 , n6201 );
or ( n7054 , n7049 , n7053 );
and ( n7055 , n7054 , n5188 );
and ( n7056 , n3776 , n5282 );
or ( n7057 , n7055 , n7056 );
and ( n7058 , n7057 , n6218 );
not ( n7059 , n6694 );
and ( n7060 , n7059 , n6356 );
xor ( n7061 , n6356 , n6345 );
and ( n7062 , n6697 , n6345 );
xor ( n7063 , n7061 , n7062 );
and ( n7064 , n7063 , n6694 );
or ( n7065 , n7060 , n7064 );
and ( n7066 , n7065 , n5188 );
and ( n7067 , n3776 , n5282 );
or ( n7068 , n7066 , n7067 );
and ( n7069 , n7068 , n6710 );
and ( n7070 , n5757 , n5188 );
and ( n7071 , n3776 , n5282 );
or ( n7072 , n7070 , n7071 );
and ( n7073 , n7072 , n6717 );
and ( n7074 , n5757 , n6719 );
not ( n7075 , n5757 );
not ( n7076 , n5492 );
xor ( n7077 , n7075 , n7076 );
and ( n7078 , n7077 , n5188 );
and ( n7079 , n3776 , n5282 );
or ( n7080 , n7078 , n7079 );
and ( n7081 , n7080 , n6724 );
or ( n7082 , n6738 , n7047 , n7058 , n7069 , n7073 , n7074 , n7081 );
and ( n7083 , n6737 , n7082 );
and ( n7084 , n3776 , n3260 );
or ( n7085 , n7083 , n7084 );
and ( n7086 , n7085 , n2422 );
and ( n7087 , n3772 , n2428 );
or ( n7088 , n7086 , n7087 );
buf ( n7089 , n7088 );
buf ( n7090 , n2424 );
buf ( n7091 , n2281 );
buf ( n7092 , n2280 );
not ( n7093 , n3260 );
and ( n7094 , n4249 , n3631 );
not ( n7095 , n7021 );
and ( n7096 , n7095 , n6749 );
xor ( n7097 , n6749 , n3770 );
and ( n7098 , n7024 , n3770 );
xor ( n7099 , n7097 , n7098 );
and ( n7100 , n7099 , n7021 );
or ( n7101 , n7096 , n7100 );
and ( n7102 , n7101 , n5289 );
and ( n7103 , n7101 , n5287 );
not ( n7104 , n3290 );
and ( n7105 , n7104 , n4599 );
not ( n7106 , n4999 );
and ( n7107 , n7106 , n4607 );
xor ( n7108 , n4607 , n4578 );
and ( n7109 , n7034 , n7035 );
xor ( n7110 , n7108 , n7109 );
and ( n7111 , n7110 , n4999 );
or ( n7112 , n7107 , n7111 );
and ( n7113 , n7112 , n3290 );
or ( n7114 , n7105 , n7113 );
and ( n7115 , n7114 , n5152 );
and ( n7116 , n4599 , n5154 );
or ( n7117 , n7102 , n7103 , n7115 , n7116 );
and ( n7118 , n7117 , n5188 );
and ( n7119 , n4249 , n5282 );
or ( n7120 , n7118 , n7119 );
and ( n7121 , n7120 , n5285 );
not ( n7122 , n6201 );
and ( n7123 , n7122 , n5875 );
xor ( n7124 , n5875 , n5852 );
and ( n7125 , n7050 , n7051 );
xor ( n7126 , n7124 , n7125 );
and ( n7127 , n7126 , n6201 );
or ( n7128 , n7123 , n7127 );
and ( n7129 , n7128 , n5188 );
and ( n7130 , n4249 , n5282 );
or ( n7131 , n7129 , n7130 );
and ( n7132 , n7131 , n6218 );
not ( n7133 , n6694 );
and ( n7134 , n7133 , n6368 );
xor ( n7135 , n6368 , n6345 );
and ( n7136 , n7061 , n7062 );
xor ( n7137 , n7135 , n7136 );
and ( n7138 , n7137 , n6694 );
or ( n7139 , n7134 , n7138 );
and ( n7140 , n7139 , n5188 );
and ( n7141 , n4249 , n5282 );
or ( n7142 , n7140 , n7141 );
and ( n7143 , n7142 , n6710 );
and ( n7144 , n5747 , n5188 );
and ( n7145 , n4249 , n5282 );
or ( n7146 , n7144 , n7145 );
and ( n7147 , n7146 , n6717 );
and ( n7148 , n5747 , n6719 );
not ( n7149 , n5747 );
and ( n7150 , n7075 , n7076 );
xor ( n7151 , n7149 , n7150 );
and ( n7152 , n7151 , n5188 );
and ( n7153 , n4249 , n5282 );
or ( n7154 , n7152 , n7153 );
and ( n7155 , n7154 , n6724 );
or ( n7156 , n7094 , n7121 , n7132 , n7143 , n7147 , n7148 , n7155 );
and ( n7157 , n7093 , n7156 );
and ( n7158 , n4249 , n3260 );
or ( n7159 , n7157 , n7158 );
and ( n7160 , n7159 , n2422 );
and ( n7161 , n4245 , n2428 );
or ( n7162 , n7160 , n7161 );
buf ( n7163 , n7162 );
buf ( n7164 , n2424 );
buf ( n7165 , n2281 );
buf ( n7166 , n2280 );
not ( n7167 , n3260 );
and ( n7168 , n4235 , n3631 );
not ( n7169 , n7021 );
and ( n7170 , n7169 , n6759 );
xor ( n7171 , n6759 , n3770 );
and ( n7172 , n7097 , n7098 );
xor ( n7173 , n7171 , n7172 );
and ( n7174 , n7173 , n7021 );
or ( n7175 , n7170 , n7174 );
and ( n7176 , n7175 , n5289 );
and ( n7177 , n7175 , n5287 );
not ( n7178 , n3290 );
and ( n7179 , n7178 , n4614 );
not ( n7180 , n4999 );
and ( n7181 , n7180 , n4622 );
xor ( n7182 , n4622 , n4578 );
and ( n7183 , n7108 , n7109 );
xor ( n7184 , n7182 , n7183 );
and ( n7185 , n7184 , n4999 );
or ( n7186 , n7181 , n7185 );
and ( n7187 , n7186 , n3290 );
or ( n7188 , n7179 , n7187 );
and ( n7189 , n7188 , n5152 );
and ( n7190 , n4614 , n5154 );
or ( n7191 , n7176 , n7177 , n7189 , n7190 );
and ( n7192 , n7191 , n5188 );
and ( n7193 , n4235 , n5282 );
or ( n7194 , n7192 , n7193 );
and ( n7195 , n7194 , n5285 );
not ( n7196 , n6201 );
and ( n7197 , n7196 , n5887 );
xor ( n7198 , n5887 , n5852 );
and ( n7199 , n7124 , n7125 );
xor ( n7200 , n7198 , n7199 );
and ( n7201 , n7200 , n6201 );
or ( n7202 , n7197 , n7201 );
and ( n7203 , n7202 , n5188 );
and ( n7204 , n4235 , n5282 );
or ( n7205 , n7203 , n7204 );
and ( n7206 , n7205 , n6218 );
not ( n7207 , n6694 );
and ( n7208 , n7207 , n6380 );
xor ( n7209 , n6380 , n6345 );
and ( n7210 , n7135 , n7136 );
xor ( n7211 , n7209 , n7210 );
and ( n7212 , n7211 , n6694 );
or ( n7213 , n7208 , n7212 );
and ( n7214 , n7213 , n5188 );
and ( n7215 , n4235 , n5282 );
or ( n7216 , n7214 , n7215 );
and ( n7217 , n7216 , n6710 );
and ( n7218 , n5737 , n5188 );
and ( n7219 , n4235 , n5282 );
or ( n7220 , n7218 , n7219 );
and ( n7221 , n7220 , n6717 );
and ( n7222 , n5737 , n6719 );
not ( n7223 , n5737 );
and ( n7224 , n7149 , n7150 );
xor ( n7225 , n7223 , n7224 );
and ( n7226 , n7225 , n5188 );
and ( n7227 , n4235 , n5282 );
or ( n7228 , n7226 , n7227 );
and ( n7229 , n7228 , n6724 );
or ( n7230 , n7168 , n7195 , n7206 , n7217 , n7221 , n7222 , n7229 );
and ( n7231 , n7167 , n7230 );
and ( n7232 , n4235 , n3260 );
or ( n7233 , n7231 , n7232 );
and ( n7234 , n7233 , n2422 );
and ( n7235 , n3945 , n2428 );
or ( n7236 , n7234 , n7235 );
buf ( n7237 , n7236 );
buf ( n7238 , n2424 );
buf ( n7239 , n2281 );
buf ( n7240 , n2280 );
not ( n7241 , n3260 );
and ( n7242 , n4225 , n3631 );
not ( n7243 , n7021 );
and ( n7244 , n7243 , n6769 );
xor ( n7245 , n6769 , n3770 );
and ( n7246 , n7171 , n7172 );
xor ( n7247 , n7245 , n7246 );
and ( n7248 , n7247 , n7021 );
or ( n7249 , n7244 , n7248 );
and ( n7250 , n7249 , n5289 );
and ( n7251 , n7249 , n5287 );
not ( n7252 , n3290 );
and ( n7253 , n7252 , n4629 );
not ( n7254 , n4999 );
and ( n7255 , n7254 , n4637 );
xor ( n7256 , n4637 , n4578 );
and ( n7257 , n7182 , n7183 );
xor ( n7258 , n7256 , n7257 );
and ( n7259 , n7258 , n4999 );
or ( n7260 , n7255 , n7259 );
and ( n7261 , n7260 , n3290 );
or ( n7262 , n7253 , n7261 );
and ( n7263 , n7262 , n5152 );
and ( n7264 , n4629 , n5154 );
or ( n7265 , n7250 , n7251 , n7263 , n7264 );
and ( n7266 , n7265 , n5188 );
and ( n7267 , n4225 , n5282 );
or ( n7268 , n7266 , n7267 );
and ( n7269 , n7268 , n5285 );
not ( n7270 , n6201 );
and ( n7271 , n7270 , n5899 );
xor ( n7272 , n5899 , n5852 );
and ( n7273 , n7198 , n7199 );
xor ( n7274 , n7272 , n7273 );
and ( n7275 , n7274 , n6201 );
or ( n7276 , n7271 , n7275 );
and ( n7277 , n7276 , n5188 );
and ( n7278 , n4225 , n5282 );
or ( n7279 , n7277 , n7278 );
and ( n7280 , n7279 , n6218 );
not ( n7281 , n6694 );
and ( n7282 , n7281 , n6392 );
xor ( n7283 , n6392 , n6345 );
and ( n7284 , n7209 , n7210 );
xor ( n7285 , n7283 , n7284 );
and ( n7286 , n7285 , n6694 );
or ( n7287 , n7282 , n7286 );
and ( n7288 , n7287 , n5188 );
and ( n7289 , n4225 , n5282 );
or ( n7290 , n7288 , n7289 );
and ( n7291 , n7290 , n6710 );
and ( n7292 , n5727 , n5188 );
and ( n7293 , n4225 , n5282 );
or ( n7294 , n7292 , n7293 );
and ( n7295 , n7294 , n6717 );
and ( n7296 , n5727 , n6719 );
not ( n7297 , n5727 );
and ( n7298 , n7223 , n7224 );
xor ( n7299 , n7297 , n7298 );
and ( n7300 , n7299 , n5188 );
and ( n7301 , n4225 , n5282 );
or ( n7302 , n7300 , n7301 );
and ( n7303 , n7302 , n6724 );
or ( n7304 , n7242 , n7269 , n7280 , n7291 , n7295 , n7296 , n7303 );
and ( n7305 , n7241 , n7304 );
and ( n7306 , n4225 , n3260 );
or ( n7307 , n7305 , n7306 );
and ( n7308 , n7307 , n2422 );
and ( n7309 , n3940 , n2428 );
or ( n7310 , n7308 , n7309 );
buf ( n7311 , n7310 );
buf ( n7312 , n2424 );
buf ( n7313 , n2281 );
buf ( n7314 , n2280 );
not ( n7315 , n3260 );
and ( n7316 , n4215 , n3631 );
not ( n7317 , n7021 );
and ( n7318 , n7317 , n6779 );
xor ( n7319 , n6779 , n3770 );
and ( n7320 , n7245 , n7246 );
xor ( n7321 , n7319 , n7320 );
and ( n7322 , n7321 , n7021 );
or ( n7323 , n7318 , n7322 );
and ( n7324 , n7323 , n5289 );
and ( n7325 , n7323 , n5287 );
not ( n7326 , n3290 );
and ( n7327 , n7326 , n4644 );
not ( n7328 , n4999 );
and ( n7329 , n7328 , n4652 );
xor ( n7330 , n4652 , n4578 );
and ( n7331 , n7256 , n7257 );
xor ( n7332 , n7330 , n7331 );
and ( n7333 , n7332 , n4999 );
or ( n7334 , n7329 , n7333 );
and ( n7335 , n7334 , n3290 );
or ( n7336 , n7327 , n7335 );
and ( n7337 , n7336 , n5152 );
and ( n7338 , n4644 , n5154 );
or ( n7339 , n7324 , n7325 , n7337 , n7338 );
and ( n7340 , n7339 , n5188 );
and ( n7341 , n4215 , n5282 );
or ( n7342 , n7340 , n7341 );
and ( n7343 , n7342 , n5285 );
not ( n7344 , n6201 );
and ( n7345 , n7344 , n5911 );
xor ( n7346 , n5911 , n5852 );
and ( n7347 , n7272 , n7273 );
xor ( n7348 , n7346 , n7347 );
and ( n7349 , n7348 , n6201 );
or ( n7350 , n7345 , n7349 );
and ( n7351 , n7350 , n5188 );
and ( n7352 , n4215 , n5282 );
or ( n7353 , n7351 , n7352 );
and ( n7354 , n7353 , n6218 );
not ( n7355 , n6694 );
and ( n7356 , n7355 , n6404 );
xor ( n7357 , n6404 , n6345 );
and ( n7358 , n7283 , n7284 );
xor ( n7359 , n7357 , n7358 );
and ( n7360 , n7359 , n6694 );
or ( n7361 , n7356 , n7360 );
and ( n7362 , n7361 , n5188 );
and ( n7363 , n4215 , n5282 );
or ( n7364 , n7362 , n7363 );
and ( n7365 , n7364 , n6710 );
and ( n7366 , n5717 , n5188 );
and ( n7367 , n4215 , n5282 );
or ( n7368 , n7366 , n7367 );
and ( n7369 , n7368 , n6717 );
and ( n7370 , n5717 , n6719 );
not ( n7371 , n5717 );
and ( n7372 , n7297 , n7298 );
xor ( n7373 , n7371 , n7372 );
and ( n7374 , n7373 , n5188 );
and ( n7375 , n4215 , n5282 );
or ( n7376 , n7374 , n7375 );
and ( n7377 , n7376 , n6724 );
or ( n7378 , n7316 , n7343 , n7354 , n7365 , n7369 , n7370 , n7377 );
and ( n7379 , n7315 , n7378 );
and ( n7380 , n4215 , n3260 );
or ( n7381 , n7379 , n7380 );
and ( n7382 , n7381 , n2422 );
and ( n7383 , n3935 , n2428 );
or ( n7384 , n7382 , n7383 );
buf ( n7385 , n7384 );
buf ( n7386 , n2424 );
buf ( n7387 , n2281 );
buf ( n7388 , n2280 );
not ( n7389 , n3260 );
and ( n7390 , n4205 , n3631 );
not ( n7391 , n7021 );
and ( n7392 , n7391 , n6789 );
xor ( n7393 , n6789 , n3770 );
and ( n7394 , n7319 , n7320 );
xor ( n7395 , n7393 , n7394 );
and ( n7396 , n7395 , n7021 );
or ( n7397 , n7392 , n7396 );
and ( n7398 , n7397 , n5289 );
and ( n7399 , n7397 , n5287 );
not ( n7400 , n3290 );
and ( n7401 , n7400 , n4659 );
not ( n7402 , n4999 );
and ( n7403 , n7402 , n4667 );
xor ( n7404 , n4667 , n4578 );
and ( n7405 , n7330 , n7331 );
xor ( n7406 , n7404 , n7405 );
and ( n7407 , n7406 , n4999 );
or ( n7408 , n7403 , n7407 );
and ( n7409 , n7408 , n3290 );
or ( n7410 , n7401 , n7409 );
and ( n7411 , n7410 , n5152 );
and ( n7412 , n4659 , n5154 );
or ( n7413 , n7398 , n7399 , n7411 , n7412 );
and ( n7414 , n7413 , n5188 );
and ( n7415 , n4205 , n5282 );
or ( n7416 , n7414 , n7415 );
and ( n7417 , n7416 , n5285 );
not ( n7418 , n6201 );
and ( n7419 , n7418 , n5923 );
xor ( n7420 , n5923 , n5852 );
and ( n7421 , n7346 , n7347 );
xor ( n7422 , n7420 , n7421 );
and ( n7423 , n7422 , n6201 );
or ( n7424 , n7419 , n7423 );
and ( n7425 , n7424 , n5188 );
and ( n7426 , n4205 , n5282 );
or ( n7427 , n7425 , n7426 );
and ( n7428 , n7427 , n6218 );
not ( n7429 , n6694 );
and ( n7430 , n7429 , n6416 );
xor ( n7431 , n6416 , n6345 );
and ( n7432 , n7357 , n7358 );
xor ( n7433 , n7431 , n7432 );
and ( n7434 , n7433 , n6694 );
or ( n7435 , n7430 , n7434 );
and ( n7436 , n7435 , n5188 );
and ( n7437 , n4205 , n5282 );
or ( n7438 , n7436 , n7437 );
and ( n7439 , n7438 , n6710 );
and ( n7440 , n5707 , n5188 );
and ( n7441 , n4205 , n5282 );
or ( n7442 , n7440 , n7441 );
and ( n7443 , n7442 , n6717 );
and ( n7444 , n5707 , n6719 );
not ( n7445 , n5707 );
and ( n7446 , n7371 , n7372 );
xor ( n7447 , n7445 , n7446 );
and ( n7448 , n7447 , n5188 );
and ( n7449 , n4205 , n5282 );
or ( n7450 , n7448 , n7449 );
and ( n7451 , n7450 , n6724 );
or ( n7452 , n7390 , n7417 , n7428 , n7439 , n7443 , n7444 , n7451 );
and ( n7453 , n7389 , n7452 );
and ( n7454 , n4205 , n3260 );
or ( n7455 , n7453 , n7454 );
and ( n7456 , n7455 , n2422 );
and ( n7457 , n3930 , n2428 );
or ( n7458 , n7456 , n7457 );
buf ( n7459 , n7458 );
buf ( n7460 , n2424 );
buf ( n7461 , n2281 );
buf ( n7462 , n2280 );
not ( n7463 , n3260 );
and ( n7464 , n4195 , n3631 );
not ( n7465 , n7021 );
and ( n7466 , n7465 , n6799 );
xor ( n7467 , n6799 , n3770 );
and ( n7468 , n7393 , n7394 );
xor ( n7469 , n7467 , n7468 );
and ( n7470 , n7469 , n7021 );
or ( n7471 , n7466 , n7470 );
and ( n7472 , n7471 , n5289 );
and ( n7473 , n7471 , n5287 );
not ( n7474 , n3290 );
and ( n7475 , n7474 , n4674 );
not ( n7476 , n4999 );
and ( n7477 , n7476 , n4682 );
xor ( n7478 , n4682 , n4578 );
and ( n7479 , n7404 , n7405 );
xor ( n7480 , n7478 , n7479 );
and ( n7481 , n7480 , n4999 );
or ( n7482 , n7477 , n7481 );
and ( n7483 , n7482 , n3290 );
or ( n7484 , n7475 , n7483 );
and ( n7485 , n7484 , n5152 );
and ( n7486 , n4674 , n5154 );
or ( n7487 , n7472 , n7473 , n7485 , n7486 );
and ( n7488 , n7487 , n5188 );
and ( n7489 , n4195 , n5282 );
or ( n7490 , n7488 , n7489 );
and ( n7491 , n7490 , n5285 );
not ( n7492 , n6201 );
and ( n7493 , n7492 , n5935 );
xor ( n7494 , n5935 , n5852 );
and ( n7495 , n7420 , n7421 );
xor ( n7496 , n7494 , n7495 );
and ( n7497 , n7496 , n6201 );
or ( n7498 , n7493 , n7497 );
and ( n7499 , n7498 , n5188 );
and ( n7500 , n4195 , n5282 );
or ( n7501 , n7499 , n7500 );
and ( n7502 , n7501 , n6218 );
not ( n7503 , n6694 );
and ( n7504 , n7503 , n6428 );
xor ( n7505 , n6428 , n6345 );
and ( n7506 , n7431 , n7432 );
xor ( n7507 , n7505 , n7506 );
and ( n7508 , n7507 , n6694 );
or ( n7509 , n7504 , n7508 );
and ( n7510 , n7509 , n5188 );
and ( n7511 , n4195 , n5282 );
or ( n7512 , n7510 , n7511 );
and ( n7513 , n7512 , n6710 );
and ( n7514 , n5697 , n5188 );
and ( n7515 , n4195 , n5282 );
or ( n7516 , n7514 , n7515 );
and ( n7517 , n7516 , n6717 );
and ( n7518 , n5697 , n6719 );
not ( n7519 , n5697 );
and ( n7520 , n7445 , n7446 );
xor ( n7521 , n7519 , n7520 );
and ( n7522 , n7521 , n5188 );
and ( n7523 , n4195 , n5282 );
or ( n7524 , n7522 , n7523 );
and ( n7525 , n7524 , n6724 );
or ( n7526 , n7464 , n7491 , n7502 , n7513 , n7517 , n7518 , n7525 );
and ( n7527 , n7463 , n7526 );
and ( n7528 , n4195 , n3260 );
or ( n7529 , n7527 , n7528 );
and ( n7530 , n7529 , n2422 );
and ( n7531 , n3925 , n2428 );
or ( n7532 , n7530 , n7531 );
buf ( n7533 , n7532 );
buf ( n7534 , n2424 );
buf ( n7535 , n2281 );
buf ( n7536 , n2280 );
not ( n7537 , n3260 );
and ( n7538 , n4185 , n3631 );
not ( n7539 , n7021 );
and ( n7540 , n7539 , n6809 );
xor ( n7541 , n6809 , n3770 );
and ( n7542 , n7467 , n7468 );
xor ( n7543 , n7541 , n7542 );
and ( n7544 , n7543 , n7021 );
or ( n7545 , n7540 , n7544 );
and ( n7546 , n7545 , n5289 );
and ( n7547 , n7545 , n5287 );
not ( n7548 , n3290 );
and ( n7549 , n7548 , n4689 );
not ( n7550 , n4999 );
and ( n7551 , n7550 , n4697 );
xor ( n7552 , n4697 , n4578 );
and ( n7553 , n7478 , n7479 );
xor ( n7554 , n7552 , n7553 );
and ( n7555 , n7554 , n4999 );
or ( n7556 , n7551 , n7555 );
and ( n7557 , n7556 , n3290 );
or ( n7558 , n7549 , n7557 );
and ( n7559 , n7558 , n5152 );
and ( n7560 , n4689 , n5154 );
or ( n7561 , n7546 , n7547 , n7559 , n7560 );
and ( n7562 , n7561 , n5188 );
and ( n7563 , n4185 , n5282 );
or ( n7564 , n7562 , n7563 );
and ( n7565 , n7564 , n5285 );
not ( n7566 , n6201 );
and ( n7567 , n7566 , n5947 );
xor ( n7568 , n5947 , n5852 );
and ( n7569 , n7494 , n7495 );
xor ( n7570 , n7568 , n7569 );
and ( n7571 , n7570 , n6201 );
or ( n7572 , n7567 , n7571 );
and ( n7573 , n7572 , n5188 );
and ( n7574 , n4185 , n5282 );
or ( n7575 , n7573 , n7574 );
and ( n7576 , n7575 , n6218 );
not ( n7577 , n6694 );
and ( n7578 , n7577 , n6440 );
xor ( n7579 , n6440 , n6345 );
and ( n7580 , n7505 , n7506 );
xor ( n7581 , n7579 , n7580 );
and ( n7582 , n7581 , n6694 );
or ( n7583 , n7578 , n7582 );
and ( n7584 , n7583 , n5188 );
and ( n7585 , n4185 , n5282 );
or ( n7586 , n7584 , n7585 );
and ( n7587 , n7586 , n6710 );
and ( n7588 , n5687 , n5188 );
and ( n7589 , n4185 , n5282 );
or ( n7590 , n7588 , n7589 );
and ( n7591 , n7590 , n6717 );
and ( n7592 , n5687 , n6719 );
not ( n7593 , n5687 );
and ( n7594 , n7519 , n7520 );
xor ( n7595 , n7593 , n7594 );
and ( n7596 , n7595 , n5188 );
and ( n7597 , n4185 , n5282 );
or ( n7598 , n7596 , n7597 );
and ( n7599 , n7598 , n6724 );
or ( n7600 , n7538 , n7565 , n7576 , n7587 , n7591 , n7592 , n7599 );
and ( n7601 , n7537 , n7600 );
and ( n7602 , n4185 , n3260 );
or ( n7603 , n7601 , n7602 );
and ( n7604 , n7603 , n2422 );
and ( n7605 , n3920 , n2428 );
or ( n7606 , n7604 , n7605 );
buf ( n7607 , n7606 );
buf ( n7608 , n2424 );
buf ( n7609 , n2281 );
buf ( n7610 , n2280 );
not ( n7611 , n3260 );
and ( n7612 , n4175 , n3631 );
not ( n7613 , n7021 );
and ( n7614 , n7613 , n6819 );
xor ( n7615 , n6819 , n3770 );
and ( n7616 , n7541 , n7542 );
xor ( n7617 , n7615 , n7616 );
and ( n7618 , n7617 , n7021 );
or ( n7619 , n7614 , n7618 );
and ( n7620 , n7619 , n5289 );
and ( n7621 , n7619 , n5287 );
not ( n7622 , n3290 );
and ( n7623 , n7622 , n4704 );
not ( n7624 , n4999 );
and ( n7625 , n7624 , n4712 );
xor ( n7626 , n4712 , n4578 );
and ( n7627 , n7552 , n7553 );
xor ( n7628 , n7626 , n7627 );
and ( n7629 , n7628 , n4999 );
or ( n7630 , n7625 , n7629 );
and ( n7631 , n7630 , n3290 );
or ( n7632 , n7623 , n7631 );
and ( n7633 , n7632 , n5152 );
and ( n7634 , n4704 , n5154 );
or ( n7635 , n7620 , n7621 , n7633 , n7634 );
and ( n7636 , n7635 , n5188 );
and ( n7637 , n4175 , n5282 );
or ( n7638 , n7636 , n7637 );
and ( n7639 , n7638 , n5285 );
not ( n7640 , n6201 );
and ( n7641 , n7640 , n5959 );
xor ( n7642 , n5959 , n5852 );
and ( n7643 , n7568 , n7569 );
xor ( n7644 , n7642 , n7643 );
and ( n7645 , n7644 , n6201 );
or ( n7646 , n7641 , n7645 );
and ( n7647 , n7646 , n5188 );
and ( n7648 , n4175 , n5282 );
or ( n7649 , n7647 , n7648 );
and ( n7650 , n7649 , n6218 );
not ( n7651 , n6694 );
and ( n7652 , n7651 , n6452 );
xor ( n7653 , n6452 , n6345 );
and ( n7654 , n7579 , n7580 );
xor ( n7655 , n7653 , n7654 );
and ( n7656 , n7655 , n6694 );
or ( n7657 , n7652 , n7656 );
and ( n7658 , n7657 , n5188 );
and ( n7659 , n4175 , n5282 );
or ( n7660 , n7658 , n7659 );
and ( n7661 , n7660 , n6710 );
and ( n7662 , n5677 , n5188 );
and ( n7663 , n4175 , n5282 );
or ( n7664 , n7662 , n7663 );
and ( n7665 , n7664 , n6717 );
and ( n7666 , n5677 , n6719 );
not ( n7667 , n5677 );
and ( n7668 , n7593 , n7594 );
xor ( n7669 , n7667 , n7668 );
and ( n7670 , n7669 , n5188 );
and ( n7671 , n4175 , n5282 );
or ( n7672 , n7670 , n7671 );
and ( n7673 , n7672 , n6724 );
or ( n7674 , n7612 , n7639 , n7650 , n7661 , n7665 , n7666 , n7673 );
and ( n7675 , n7611 , n7674 );
and ( n7676 , n4175 , n3260 );
or ( n7677 , n7675 , n7676 );
and ( n7678 , n7677 , n2422 );
and ( n7679 , n3915 , n2428 );
or ( n7680 , n7678 , n7679 );
buf ( n7681 , n7680 );
buf ( n7682 , n2424 );
buf ( n7683 , n2281 );
buf ( n7684 , n2280 );
not ( n7685 , n3260 );
and ( n7686 , n4165 , n3631 );
not ( n7687 , n7021 );
and ( n7688 , n7687 , n6829 );
xor ( n7689 , n6829 , n3770 );
and ( n7690 , n7615 , n7616 );
xor ( n7691 , n7689 , n7690 );
and ( n7692 , n7691 , n7021 );
or ( n7693 , n7688 , n7692 );
and ( n7694 , n7693 , n5289 );
and ( n7695 , n7693 , n5287 );
not ( n7696 , n3290 );
and ( n7697 , n7696 , n4719 );
not ( n7698 , n4999 );
and ( n7699 , n7698 , n4727 );
xor ( n7700 , n4727 , n4578 );
and ( n7701 , n7626 , n7627 );
xor ( n7702 , n7700 , n7701 );
and ( n7703 , n7702 , n4999 );
or ( n7704 , n7699 , n7703 );
and ( n7705 , n7704 , n3290 );
or ( n7706 , n7697 , n7705 );
and ( n7707 , n7706 , n5152 );
and ( n7708 , n4719 , n5154 );
or ( n7709 , n7694 , n7695 , n7707 , n7708 );
and ( n7710 , n7709 , n5188 );
and ( n7711 , n4165 , n5282 );
or ( n7712 , n7710 , n7711 );
and ( n7713 , n7712 , n5285 );
not ( n7714 , n6201 );
and ( n7715 , n7714 , n5971 );
xor ( n7716 , n5971 , n5852 );
and ( n7717 , n7642 , n7643 );
xor ( n7718 , n7716 , n7717 );
and ( n7719 , n7718 , n6201 );
or ( n7720 , n7715 , n7719 );
and ( n7721 , n7720 , n5188 );
and ( n7722 , n4165 , n5282 );
or ( n7723 , n7721 , n7722 );
and ( n7724 , n7723 , n6218 );
not ( n7725 , n6694 );
and ( n7726 , n7725 , n6464 );
xor ( n7727 , n6464 , n6345 );
and ( n7728 , n7653 , n7654 );
xor ( n7729 , n7727 , n7728 );
and ( n7730 , n7729 , n6694 );
or ( n7731 , n7726 , n7730 );
and ( n7732 , n7731 , n5188 );
and ( n7733 , n4165 , n5282 );
or ( n7734 , n7732 , n7733 );
and ( n7735 , n7734 , n6710 );
and ( n7736 , n5667 , n5188 );
and ( n7737 , n4165 , n5282 );
or ( n7738 , n7736 , n7737 );
and ( n7739 , n7738 , n6717 );
and ( n7740 , n5667 , n6719 );
not ( n7741 , n5667 );
and ( n7742 , n7667 , n7668 );
xor ( n7743 , n7741 , n7742 );
and ( n7744 , n7743 , n5188 );
and ( n7745 , n4165 , n5282 );
or ( n7746 , n7744 , n7745 );
and ( n7747 , n7746 , n6724 );
or ( n7748 , n7686 , n7713 , n7724 , n7735 , n7739 , n7740 , n7747 );
and ( n7749 , n7685 , n7748 );
and ( n7750 , n4165 , n3260 );
or ( n7751 , n7749 , n7750 );
and ( n7752 , n7751 , n2422 );
and ( n7753 , n3910 , n2428 );
or ( n7754 , n7752 , n7753 );
buf ( n7755 , n7754 );
buf ( n7756 , n2424 );
buf ( n7757 , n2281 );
buf ( n7758 , n2280 );
not ( n7759 , n3260 );
and ( n7760 , n4155 , n3631 );
not ( n7761 , n7021 );
and ( n7762 , n7761 , n6839 );
xor ( n7763 , n6839 , n3770 );
and ( n7764 , n7689 , n7690 );
xor ( n7765 , n7763 , n7764 );
and ( n7766 , n7765 , n7021 );
or ( n7767 , n7762 , n7766 );
and ( n7768 , n7767 , n5289 );
and ( n7769 , n7767 , n5287 );
not ( n7770 , n3290 );
and ( n7771 , n7770 , n4734 );
not ( n7772 , n4999 );
and ( n7773 , n7772 , n4742 );
xor ( n7774 , n4742 , n4578 );
and ( n7775 , n7700 , n7701 );
xor ( n7776 , n7774 , n7775 );
and ( n7777 , n7776 , n4999 );
or ( n7778 , n7773 , n7777 );
and ( n7779 , n7778 , n3290 );
or ( n7780 , n7771 , n7779 );
and ( n7781 , n7780 , n5152 );
and ( n7782 , n4734 , n5154 );
or ( n7783 , n7768 , n7769 , n7781 , n7782 );
and ( n7784 , n7783 , n5188 );
and ( n7785 , n4155 , n5282 );
or ( n7786 , n7784 , n7785 );
and ( n7787 , n7786 , n5285 );
not ( n7788 , n6201 );
and ( n7789 , n7788 , n5983 );
xor ( n7790 , n5983 , n5852 );
and ( n7791 , n7716 , n7717 );
xor ( n7792 , n7790 , n7791 );
and ( n7793 , n7792 , n6201 );
or ( n7794 , n7789 , n7793 );
and ( n7795 , n7794 , n5188 );
and ( n7796 , n4155 , n5282 );
or ( n7797 , n7795 , n7796 );
and ( n7798 , n7797 , n6218 );
not ( n7799 , n6694 );
and ( n7800 , n7799 , n6476 );
xor ( n7801 , n6476 , n6345 );
and ( n7802 , n7727 , n7728 );
xor ( n7803 , n7801 , n7802 );
and ( n7804 , n7803 , n6694 );
or ( n7805 , n7800 , n7804 );
and ( n7806 , n7805 , n5188 );
and ( n7807 , n4155 , n5282 );
or ( n7808 , n7806 , n7807 );
and ( n7809 , n7808 , n6710 );
and ( n7810 , n5657 , n5188 );
and ( n7811 , n4155 , n5282 );
or ( n7812 , n7810 , n7811 );
and ( n7813 , n7812 , n6717 );
and ( n7814 , n5657 , n6719 );
not ( n7815 , n5657 );
and ( n7816 , n7741 , n7742 );
xor ( n7817 , n7815 , n7816 );
and ( n7818 , n7817 , n5188 );
and ( n7819 , n4155 , n5282 );
or ( n7820 , n7818 , n7819 );
and ( n7821 , n7820 , n6724 );
or ( n7822 , n7760 , n7787 , n7798 , n7809 , n7813 , n7814 , n7821 );
and ( n7823 , n7759 , n7822 );
and ( n7824 , n4155 , n3260 );
or ( n7825 , n7823 , n7824 );
and ( n7826 , n7825 , n2422 );
and ( n7827 , n3905 , n2428 );
or ( n7828 , n7826 , n7827 );
buf ( n7829 , n7828 );
buf ( n7830 , n2424 );
buf ( n7831 , n2281 );
buf ( n7832 , n2280 );
not ( n7833 , n3260 );
and ( n7834 , n4145 , n3631 );
not ( n7835 , n7021 );
and ( n7836 , n7835 , n6849 );
xor ( n7837 , n6849 , n3770 );
and ( n7838 , n7763 , n7764 );
xor ( n7839 , n7837 , n7838 );
and ( n7840 , n7839 , n7021 );
or ( n7841 , n7836 , n7840 );
and ( n7842 , n7841 , n5289 );
and ( n7843 , n7841 , n5287 );
not ( n7844 , n3290 );
and ( n7845 , n7844 , n4749 );
not ( n7846 , n4999 );
and ( n7847 , n7846 , n4757 );
xor ( n7848 , n4757 , n4578 );
and ( n7849 , n7774 , n7775 );
xor ( n7850 , n7848 , n7849 );
and ( n7851 , n7850 , n4999 );
or ( n7852 , n7847 , n7851 );
and ( n7853 , n7852 , n3290 );
or ( n7854 , n7845 , n7853 );
and ( n7855 , n7854 , n5152 );
and ( n7856 , n4749 , n5154 );
or ( n7857 , n7842 , n7843 , n7855 , n7856 );
and ( n7858 , n7857 , n5188 );
and ( n7859 , n4145 , n5282 );
or ( n7860 , n7858 , n7859 );
and ( n7861 , n7860 , n5285 );
not ( n7862 , n6201 );
and ( n7863 , n7862 , n5995 );
xor ( n7864 , n5995 , n5852 );
and ( n7865 , n7790 , n7791 );
xor ( n7866 , n7864 , n7865 );
and ( n7867 , n7866 , n6201 );
or ( n7868 , n7863 , n7867 );
and ( n7869 , n7868 , n5188 );
and ( n7870 , n4145 , n5282 );
or ( n7871 , n7869 , n7870 );
and ( n7872 , n7871 , n6218 );
not ( n7873 , n6694 );
and ( n7874 , n7873 , n6488 );
xor ( n7875 , n6488 , n6345 );
and ( n7876 , n7801 , n7802 );
xor ( n7877 , n7875 , n7876 );
and ( n7878 , n7877 , n6694 );
or ( n7879 , n7874 , n7878 );
and ( n7880 , n7879 , n5188 );
and ( n7881 , n4145 , n5282 );
or ( n7882 , n7880 , n7881 );
and ( n7883 , n7882 , n6710 );
and ( n7884 , n5647 , n5188 );
and ( n7885 , n4145 , n5282 );
or ( n7886 , n7884 , n7885 );
and ( n7887 , n7886 , n6717 );
and ( n7888 , n5647 , n6719 );
not ( n7889 , n5647 );
and ( n7890 , n7815 , n7816 );
xor ( n7891 , n7889 , n7890 );
and ( n7892 , n7891 , n5188 );
and ( n7893 , n4145 , n5282 );
or ( n7894 , n7892 , n7893 );
and ( n7895 , n7894 , n6724 );
or ( n7896 , n7834 , n7861 , n7872 , n7883 , n7887 , n7888 , n7895 );
and ( n7897 , n7833 , n7896 );
and ( n7898 , n4145 , n3260 );
or ( n7899 , n7897 , n7898 );
and ( n7900 , n7899 , n2422 );
and ( n7901 , n3900 , n2428 );
or ( n7902 , n7900 , n7901 );
buf ( n7903 , n7902 );
buf ( n7904 , n2424 );
buf ( n7905 , n2281 );
buf ( n7906 , n2280 );
not ( n7907 , n3260 );
and ( n7908 , n4135 , n3631 );
not ( n7909 , n7021 );
and ( n7910 , n7909 , n6859 );
xor ( n7911 , n6859 , n3770 );
and ( n7912 , n7837 , n7838 );
xor ( n7913 , n7911 , n7912 );
and ( n7914 , n7913 , n7021 );
or ( n7915 , n7910 , n7914 );
and ( n7916 , n7915 , n5289 );
and ( n7917 , n7915 , n5287 );
not ( n7918 , n3290 );
and ( n7919 , n7918 , n4764 );
not ( n7920 , n4999 );
and ( n7921 , n7920 , n4772 );
xor ( n7922 , n4772 , n4578 );
and ( n7923 , n7848 , n7849 );
xor ( n7924 , n7922 , n7923 );
and ( n7925 , n7924 , n4999 );
or ( n7926 , n7921 , n7925 );
and ( n7927 , n7926 , n3290 );
or ( n7928 , n7919 , n7927 );
and ( n7929 , n7928 , n5152 );
and ( n7930 , n4764 , n5154 );
or ( n7931 , n7916 , n7917 , n7929 , n7930 );
and ( n7932 , n7931 , n5188 );
and ( n7933 , n4135 , n5282 );
or ( n7934 , n7932 , n7933 );
and ( n7935 , n7934 , n5285 );
not ( n7936 , n6201 );
and ( n7937 , n7936 , n6007 );
xor ( n7938 , n6007 , n5852 );
and ( n7939 , n7864 , n7865 );
xor ( n7940 , n7938 , n7939 );
and ( n7941 , n7940 , n6201 );
or ( n7942 , n7937 , n7941 );
and ( n7943 , n7942 , n5188 );
and ( n7944 , n4135 , n5282 );
or ( n7945 , n7943 , n7944 );
and ( n7946 , n7945 , n6218 );
not ( n7947 , n6694 );
and ( n7948 , n7947 , n6500 );
xor ( n7949 , n6500 , n6345 );
and ( n7950 , n7875 , n7876 );
xor ( n7951 , n7949 , n7950 );
and ( n7952 , n7951 , n6694 );
or ( n7953 , n7948 , n7952 );
and ( n7954 , n7953 , n5188 );
and ( n7955 , n4135 , n5282 );
or ( n7956 , n7954 , n7955 );
and ( n7957 , n7956 , n6710 );
and ( n7958 , n5637 , n5188 );
and ( n7959 , n4135 , n5282 );
or ( n7960 , n7958 , n7959 );
and ( n7961 , n7960 , n6717 );
and ( n7962 , n5637 , n6719 );
not ( n7963 , n5637 );
and ( n7964 , n7889 , n7890 );
xor ( n7965 , n7963 , n7964 );
and ( n7966 , n7965 , n5188 );
and ( n7967 , n4135 , n5282 );
or ( n7968 , n7966 , n7967 );
and ( n7969 , n7968 , n6724 );
or ( n7970 , n7908 , n7935 , n7946 , n7957 , n7961 , n7962 , n7969 );
and ( n7971 , n7907 , n7970 );
and ( n7972 , n4135 , n3260 );
or ( n7973 , n7971 , n7972 );
and ( n7974 , n7973 , n2422 );
and ( n7975 , n3895 , n2428 );
or ( n7976 , n7974 , n7975 );
buf ( n7977 , n7976 );
buf ( n7978 , n2424 );
buf ( n7979 , n2281 );
buf ( n7980 , n2280 );
not ( n7981 , n3260 );
and ( n7982 , n4125 , n3631 );
not ( n7983 , n7021 );
and ( n7984 , n7983 , n6869 );
xor ( n7985 , n6869 , n3770 );
and ( n7986 , n7911 , n7912 );
xor ( n7987 , n7985 , n7986 );
and ( n7988 , n7987 , n7021 );
or ( n7989 , n7984 , n7988 );
and ( n7990 , n7989 , n5289 );
and ( n7991 , n7989 , n5287 );
not ( n7992 , n3290 );
and ( n7993 , n7992 , n4779 );
not ( n7994 , n4999 );
and ( n7995 , n7994 , n4787 );
xor ( n7996 , n4787 , n4578 );
and ( n7997 , n7922 , n7923 );
xor ( n7998 , n7996 , n7997 );
and ( n7999 , n7998 , n4999 );
or ( n8000 , n7995 , n7999 );
and ( n8001 , n8000 , n3290 );
or ( n8002 , n7993 , n8001 );
and ( n8003 , n8002 , n5152 );
and ( n8004 , n4779 , n5154 );
or ( n8005 , n7990 , n7991 , n8003 , n8004 );
and ( n8006 , n8005 , n5188 );
and ( n8007 , n4125 , n5282 );
or ( n8008 , n8006 , n8007 );
and ( n8009 , n8008 , n5285 );
not ( n8010 , n6201 );
and ( n8011 , n8010 , n6019 );
xor ( n8012 , n6019 , n5852 );
and ( n8013 , n7938 , n7939 );
xor ( n8014 , n8012 , n8013 );
and ( n8015 , n8014 , n6201 );
or ( n8016 , n8011 , n8015 );
and ( n8017 , n8016 , n5188 );
and ( n8018 , n4125 , n5282 );
or ( n8019 , n8017 , n8018 );
and ( n8020 , n8019 , n6218 );
not ( n8021 , n6694 );
and ( n8022 , n8021 , n6512 );
xor ( n8023 , n6512 , n6345 );
and ( n8024 , n7949 , n7950 );
xor ( n8025 , n8023 , n8024 );
and ( n8026 , n8025 , n6694 );
or ( n8027 , n8022 , n8026 );
and ( n8028 , n8027 , n5188 );
and ( n8029 , n4125 , n5282 );
or ( n8030 , n8028 , n8029 );
and ( n8031 , n8030 , n6710 );
and ( n8032 , n5627 , n5188 );
and ( n8033 , n4125 , n5282 );
or ( n8034 , n8032 , n8033 );
and ( n8035 , n8034 , n6717 );
and ( n8036 , n5627 , n6719 );
not ( n8037 , n5627 );
and ( n8038 , n7963 , n7964 );
xor ( n8039 , n8037 , n8038 );
and ( n8040 , n8039 , n5188 );
and ( n8041 , n4125 , n5282 );
or ( n8042 , n8040 , n8041 );
and ( n8043 , n8042 , n6724 );
or ( n8044 , n7982 , n8009 , n8020 , n8031 , n8035 , n8036 , n8043 );
and ( n8045 , n7981 , n8044 );
and ( n8046 , n4125 , n3260 );
or ( n8047 , n8045 , n8046 );
and ( n8048 , n8047 , n2422 );
and ( n8049 , n3890 , n2428 );
or ( n8050 , n8048 , n8049 );
buf ( n8051 , n8050 );
buf ( n8052 , n2424 );
buf ( n8053 , n2281 );
buf ( n8054 , n2280 );
not ( n8055 , n3260 );
and ( n8056 , n4115 , n3631 );
not ( n8057 , n7021 );
and ( n8058 , n8057 , n6879 );
xor ( n8059 , n6879 , n3770 );
and ( n8060 , n7985 , n7986 );
xor ( n8061 , n8059 , n8060 );
and ( n8062 , n8061 , n7021 );
or ( n8063 , n8058 , n8062 );
and ( n8064 , n8063 , n5289 );
and ( n8065 , n8063 , n5287 );
not ( n8066 , n3290 );
and ( n8067 , n8066 , n4794 );
not ( n8068 , n4999 );
and ( n8069 , n8068 , n4802 );
xor ( n8070 , n4802 , n4578 );
and ( n8071 , n7996 , n7997 );
xor ( n8072 , n8070 , n8071 );
and ( n8073 , n8072 , n4999 );
or ( n8074 , n8069 , n8073 );
and ( n8075 , n8074 , n3290 );
or ( n8076 , n8067 , n8075 );
and ( n8077 , n8076 , n5152 );
and ( n8078 , n4794 , n5154 );
or ( n8079 , n8064 , n8065 , n8077 , n8078 );
and ( n8080 , n8079 , n5188 );
and ( n8081 , n4115 , n5282 );
or ( n8082 , n8080 , n8081 );
and ( n8083 , n8082 , n5285 );
not ( n8084 , n6201 );
and ( n8085 , n8084 , n6031 );
xor ( n8086 , n6031 , n5852 );
and ( n8087 , n8012 , n8013 );
xor ( n8088 , n8086 , n8087 );
and ( n8089 , n8088 , n6201 );
or ( n8090 , n8085 , n8089 );
and ( n8091 , n8090 , n5188 );
and ( n8092 , n4115 , n5282 );
or ( n8093 , n8091 , n8092 );
and ( n8094 , n8093 , n6218 );
not ( n8095 , n6694 );
and ( n8096 , n8095 , n6524 );
xor ( n8097 , n6524 , n6345 );
and ( n8098 , n8023 , n8024 );
xor ( n8099 , n8097 , n8098 );
and ( n8100 , n8099 , n6694 );
or ( n8101 , n8096 , n8100 );
and ( n8102 , n8101 , n5188 );
and ( n8103 , n4115 , n5282 );
or ( n8104 , n8102 , n8103 );
and ( n8105 , n8104 , n6710 );
and ( n8106 , n5617 , n5188 );
and ( n8107 , n4115 , n5282 );
or ( n8108 , n8106 , n8107 );
and ( n8109 , n8108 , n6717 );
and ( n8110 , n5617 , n6719 );
not ( n8111 , n5617 );
and ( n8112 , n8037 , n8038 );
xor ( n8113 , n8111 , n8112 );
and ( n8114 , n8113 , n5188 );
and ( n8115 , n4115 , n5282 );
or ( n8116 , n8114 , n8115 );
and ( n8117 , n8116 , n6724 );
or ( n8118 , n8056 , n8083 , n8094 , n8105 , n8109 , n8110 , n8117 );
and ( n8119 , n8055 , n8118 );
and ( n8120 , n4115 , n3260 );
or ( n8121 , n8119 , n8120 );
and ( n8122 , n8121 , n2422 );
and ( n8123 , n3885 , n2428 );
or ( n8124 , n8122 , n8123 );
buf ( n8125 , n8124 );
buf ( n8126 , n2424 );
buf ( n8127 , n2281 );
buf ( n8128 , n2280 );
not ( n8129 , n3260 );
and ( n8130 , n4105 , n3631 );
not ( n8131 , n7021 );
and ( n8132 , n8131 , n6889 );
xor ( n8133 , n6889 , n3770 );
and ( n8134 , n8059 , n8060 );
xor ( n8135 , n8133 , n8134 );
and ( n8136 , n8135 , n7021 );
or ( n8137 , n8132 , n8136 );
and ( n8138 , n8137 , n5289 );
and ( n8139 , n8137 , n5287 );
not ( n8140 , n3290 );
and ( n8141 , n8140 , n4809 );
not ( n8142 , n4999 );
and ( n8143 , n8142 , n4817 );
xor ( n8144 , n4817 , n4578 );
and ( n8145 , n8070 , n8071 );
xor ( n8146 , n8144 , n8145 );
and ( n8147 , n8146 , n4999 );
or ( n8148 , n8143 , n8147 );
and ( n8149 , n8148 , n3290 );
or ( n8150 , n8141 , n8149 );
and ( n8151 , n8150 , n5152 );
and ( n8152 , n4809 , n5154 );
or ( n8153 , n8138 , n8139 , n8151 , n8152 );
and ( n8154 , n8153 , n5188 );
and ( n8155 , n4105 , n5282 );
or ( n8156 , n8154 , n8155 );
and ( n8157 , n8156 , n5285 );
not ( n8158 , n6201 );
and ( n8159 , n8158 , n6043 );
xor ( n8160 , n6043 , n5852 );
and ( n8161 , n8086 , n8087 );
xor ( n8162 , n8160 , n8161 );
and ( n8163 , n8162 , n6201 );
or ( n8164 , n8159 , n8163 );
and ( n8165 , n8164 , n5188 );
and ( n8166 , n4105 , n5282 );
or ( n8167 , n8165 , n8166 );
and ( n8168 , n8167 , n6218 );
not ( n8169 , n6694 );
and ( n8170 , n8169 , n6536 );
xor ( n8171 , n6536 , n6345 );
and ( n8172 , n8097 , n8098 );
xor ( n8173 , n8171 , n8172 );
and ( n8174 , n8173 , n6694 );
or ( n8175 , n8170 , n8174 );
and ( n8176 , n8175 , n5188 );
and ( n8177 , n4105 , n5282 );
or ( n8178 , n8176 , n8177 );
and ( n8179 , n8178 , n6710 );
and ( n8180 , n5607 , n5188 );
and ( n8181 , n4105 , n5282 );
or ( n8182 , n8180 , n8181 );
and ( n8183 , n8182 , n6717 );
and ( n8184 , n5607 , n6719 );
not ( n8185 , n5607 );
and ( n8186 , n8111 , n8112 );
xor ( n8187 , n8185 , n8186 );
and ( n8188 , n8187 , n5188 );
and ( n8189 , n4105 , n5282 );
or ( n8190 , n8188 , n8189 );
and ( n8191 , n8190 , n6724 );
or ( n8192 , n8130 , n8157 , n8168 , n8179 , n8183 , n8184 , n8191 );
and ( n8193 , n8129 , n8192 );
and ( n8194 , n4105 , n3260 );
or ( n8195 , n8193 , n8194 );
and ( n8196 , n8195 , n2422 );
and ( n8197 , n3880 , n2428 );
or ( n8198 , n8196 , n8197 );
buf ( n8199 , n8198 );
buf ( n8200 , n2424 );
buf ( n8201 , n2281 );
buf ( n8202 , n2280 );
not ( n8203 , n3260 );
and ( n8204 , n4095 , n3631 );
not ( n8205 , n7021 );
and ( n8206 , n8205 , n6899 );
xor ( n8207 , n6899 , n3770 );
and ( n8208 , n8133 , n8134 );
xor ( n8209 , n8207 , n8208 );
and ( n8210 , n8209 , n7021 );
or ( n8211 , n8206 , n8210 );
and ( n8212 , n8211 , n5289 );
and ( n8213 , n8211 , n5287 );
not ( n8214 , n3290 );
and ( n8215 , n8214 , n4824 );
not ( n8216 , n4999 );
and ( n8217 , n8216 , n4832 );
xor ( n8218 , n4832 , n4578 );
and ( n8219 , n8144 , n8145 );
xor ( n8220 , n8218 , n8219 );
and ( n8221 , n8220 , n4999 );
or ( n8222 , n8217 , n8221 );
and ( n8223 , n8222 , n3290 );
or ( n8224 , n8215 , n8223 );
and ( n8225 , n8224 , n5152 );
and ( n8226 , n4824 , n5154 );
or ( n8227 , n8212 , n8213 , n8225 , n8226 );
and ( n8228 , n8227 , n5188 );
and ( n8229 , n4095 , n5282 );
nor ( n8230 , n8228 , n8229 );
and ( n8231 , n8230 , n5285 );
not ( n8232 , n6201 );
and ( n8233 , n8232 , n6055 );
xor ( n8234 , n6055 , n5852 );
and ( n8235 , n8160 , n8161 );
xor ( n8236 , n8234 , n8235 );
and ( n8237 , n8236 , n6201 );
or ( n8238 , n8233 , n8237 );
and ( n8239 , n8238 , n5188 );
and ( n8240 , n4095 , n5282 );
or ( n8241 , n8239 , n8240 );
and ( n8242 , n8241 , n6218 );
not ( n8243 , n6694 );
and ( n8244 , n8243 , n6548 );
xor ( n8245 , n6548 , n6345 );
and ( n8246 , n8171 , n8172 );
xor ( n8247 , n8245 , n8246 );
and ( n8248 , n8247 , n6694 );
or ( n8249 , n8244 , n8248 );
and ( n8250 , n8249 , n5188 );
and ( n8251 , n4095 , n5282 );
or ( n8252 , n8250 , n8251 );
and ( n8253 , n8252 , n6710 );
and ( n8254 , n5597 , n5188 );
and ( n8255 , n4095 , n5282 );
or ( n8256 , n8254 , n8255 );
and ( n8257 , n8256 , n6717 );
and ( n8258 , n5597 , n6719 );
not ( n8259 , n5597 );
and ( n8260 , n8185 , n8186 );
xor ( n8261 , n8259 , n8260 );
and ( n8262 , n8261 , n5188 );
and ( n8263 , n4095 , n5282 );
or ( n8264 , n8262 , n8263 );
and ( n8265 , n8264 , n6724 );
or ( n8266 , n8204 , n8231 , n8242 , n8253 , n8257 , n8258 , n8265 );
and ( n8267 , n8203 , n8266 );
and ( n8268 , n4095 , n3260 );
or ( n8269 , n8267 , n8268 );
and ( n8270 , n8269 , n2422 );
and ( n8271 , n3875 , n2428 );
or ( n8272 , n8270 , n8271 );
buf ( n8273 , n8272 );
buf ( n8274 , n2424 );
buf ( n8275 , n2281 );
buf ( n8276 , n2280 );
not ( n8277 , n3260 );
and ( n8278 , n4085 , n3631 );
not ( n8279 , n7021 );
and ( n8280 , n8279 , n6909 );
xor ( n8281 , n6909 , n3770 );
and ( n8282 , n8207 , n8208 );
xor ( n8283 , n8281 , n8282 );
and ( n8284 , n8283 , n7021 );
or ( n8285 , n8280 , n8284 );
and ( n8286 , n8285 , n5289 );
and ( n8287 , n8285 , n5287 );
not ( n8288 , n3290 );
and ( n8289 , n8288 , n4839 );
not ( n8290 , n4999 );
and ( n8291 , n8290 , n4847 );
xor ( n8292 , n4847 , n4578 );
and ( n8293 , n8218 , n8219 );
xor ( n8294 , n8292 , n8293 );
and ( n8295 , n8294 , n4999 );
or ( n8296 , n8291 , n8295 );
and ( n8297 , n8296 , n3290 );
or ( n8298 , n8289 , n8297 );
and ( n8299 , n8298 , n5152 );
and ( n8300 , n4839 , n5154 );
or ( n8301 , n8286 , n8287 , n8299 , n8300 );
and ( n8302 , n8301 , n5188 );
and ( n8303 , n4085 , n5282 );
or ( n8304 , n8302 , n8303 );
and ( n8305 , n8304 , n5285 );
not ( n8306 , n6201 );
and ( n8307 , n8306 , n6067 );
xor ( n8308 , n6067 , n5852 );
and ( n8309 , n8234 , n8235 );
xor ( n8310 , n8308 , n8309 );
and ( n8311 , n8310 , n6201 );
or ( n8312 , n8307 , n8311 );
and ( n8313 , n8312 , n5188 );
and ( n8314 , n4085 , n5282 );
or ( n8315 , n8313 , n8314 );
and ( n8316 , n8315 , n6218 );
not ( n8317 , n6694 );
and ( n8318 , n8317 , n6560 );
xor ( n8319 , n6560 , n6345 );
and ( n8320 , n8245 , n8246 );
xor ( n8321 , n8319 , n8320 );
and ( n8322 , n8321 , n6694 );
or ( n8323 , n8318 , n8322 );
and ( n8324 , n8323 , n5188 );
and ( n8325 , n4085 , n5282 );
or ( n8326 , n8324 , n8325 );
and ( n8327 , n8326 , n6710 );
and ( n8328 , n5587 , n5188 );
and ( n8329 , n4085 , n5282 );
or ( n8330 , n8328 , n8329 );
and ( n8331 , n8330 , n6717 );
and ( n8332 , n5587 , n6719 );
not ( n8333 , n5587 );
and ( n8334 , n8259 , n8260 );
xor ( n8335 , n8333 , n8334 );
and ( n8336 , n8335 , n5188 );
and ( n8337 , n4085 , n5282 );
or ( n8338 , n8336 , n8337 );
and ( n8339 , n8338 , n6724 );
or ( n8340 , n8278 , n8305 , n8316 , n8327 , n8331 , n8332 , n8339 );
and ( n8341 , n8277 , n8340 );
and ( n8342 , n4085 , n3260 );
or ( n8343 , n8341 , n8342 );
and ( n8344 , n8343 , n2422 );
and ( n8345 , n3870 , n2428 );
or ( n8346 , n8344 , n8345 );
buf ( n8347 , n8346 );
buf ( n8348 , n2424 );
buf ( n8349 , n2281 );
buf ( n8350 , n2280 );
not ( n8351 , n3260 );
and ( n8352 , n4075 , n3631 );
not ( n8353 , n7021 );
and ( n8354 , n8353 , n6919 );
xor ( n8355 , n6919 , n3770 );
and ( n8356 , n8281 , n8282 );
xor ( n8357 , n8355 , n8356 );
and ( n8358 , n8357 , n7021 );
or ( n8359 , n8354 , n8358 );
and ( n8360 , n8359 , n5289 );
and ( n8361 , n8359 , n5287 );
not ( n8362 , n3290 );
and ( n8363 , n8362 , n4854 );
not ( n8364 , n4999 );
and ( n8365 , n8364 , n4862 );
xor ( n8366 , n4862 , n4578 );
and ( n8367 , n8292 , n8293 );
xor ( n8368 , n8366 , n8367 );
and ( n8369 , n8368 , n4999 );
or ( n8370 , n8365 , n8369 );
and ( n8371 , n8370 , n3290 );
or ( n8372 , n8363 , n8371 );
and ( n8373 , n8372 , n5152 );
and ( n8374 , n4854 , n5154 );
or ( n8375 , n8360 , n8361 , n8373 , n8374 );
and ( n8376 , n8375 , n5188 );
and ( n8377 , n4075 , n5282 );
or ( n8378 , n8376 , n8377 );
and ( n8379 , n8378 , n5285 );
not ( n8380 , n6201 );
and ( n8381 , n8380 , n6079 );
xor ( n8382 , n6079 , n5852 );
and ( n8383 , n8308 , n8309 );
xor ( n8384 , n8382 , n8383 );
and ( n8385 , n8384 , n6201 );
or ( n8386 , n8381 , n8385 );
and ( n8387 , n8386 , n5188 );
and ( n8388 , n4075 , n5282 );
or ( n8389 , n8387 , n8388 );
and ( n8390 , n8389 , n6218 );
not ( n8391 , n6694 );
and ( n8392 , n8391 , n6572 );
xor ( n8393 , n6572 , n6345 );
and ( n8394 , n8319 , n8320 );
xor ( n8395 , n8393 , n8394 );
and ( n8396 , n8395 , n6694 );
or ( n8397 , n8392 , n8396 );
and ( n8398 , n8397 , n5188 );
and ( n8399 , n4075 , n5282 );
or ( n8400 , n8398 , n8399 );
and ( n8401 , n8400 , n6710 );
and ( n8402 , n5577 , n5188 );
and ( n8403 , n4075 , n5282 );
or ( n8404 , n8402 , n8403 );
and ( n8405 , n8404 , n6717 );
and ( n8406 , n5577 , n6719 );
not ( n8407 , n5577 );
and ( n8408 , n8333 , n8334 );
xor ( n8409 , n8407 , n8408 );
and ( n8410 , n8409 , n5188 );
and ( n8411 , n4075 , n5282 );
or ( n8412 , n8410 , n8411 );
and ( n8413 , n8412 , n6724 );
or ( n8414 , n8352 , n8379 , n8390 , n8401 , n8405 , n8406 , n8413 );
and ( n8415 , n8351 , n8414 );
and ( n8416 , n4075 , n3260 );
or ( n8417 , n8415 , n8416 );
and ( n8418 , n8417 , n2422 );
and ( n8419 , n3865 , n2428 );
or ( n8420 , n8418 , n8419 );
buf ( n8421 , n8420 );
buf ( n8422 , n2424 );
buf ( n8423 , n2281 );
buf ( n8424 , n2280 );
not ( n8425 , n3260 );
and ( n8426 , n4065 , n3631 );
not ( n8427 , n7021 );
and ( n8428 , n8427 , n6929 );
xor ( n8429 , n6929 , n3770 );
and ( n8430 , n8355 , n8356 );
xor ( n8431 , n8429 , n8430 );
and ( n8432 , n8431 , n7021 );
or ( n8433 , n8428 , n8432 );
and ( n8434 , n8433 , n5289 );
and ( n8435 , n8433 , n5287 );
not ( n8436 , n3290 );
and ( n8437 , n8436 , n4869 );
not ( n8438 , n4999 );
and ( n8439 , n8438 , n4877 );
xor ( n8440 , n4877 , n4578 );
and ( n8441 , n8366 , n8367 );
xor ( n8442 , n8440 , n8441 );
and ( n8443 , n8442 , n4999 );
or ( n8444 , n8439 , n8443 );
and ( n8445 , n8444 , n3290 );
or ( n8446 , n8437 , n8445 );
and ( n8447 , n8446 , n5152 );
and ( n8448 , n4869 , n5154 );
or ( n8449 , n8434 , n8435 , n8447 , n8448 );
and ( n8450 , n8449 , n5188 );
and ( n8451 , n4065 , n5282 );
or ( n8452 , n8450 , n8451 );
and ( n8453 , n8452 , n5285 );
not ( n8454 , n6201 );
and ( n8455 , n8454 , n6091 );
xor ( n8456 , n6091 , n5852 );
and ( n8457 , n8382 , n8383 );
xor ( n8458 , n8456 , n8457 );
and ( n8459 , n8458 , n6201 );
or ( n8460 , n8455 , n8459 );
and ( n8461 , n8460 , n5188 );
and ( n8462 , n4065 , n5282 );
or ( n8463 , n8461 , n8462 );
and ( n8464 , n8463 , n6218 );
not ( n8465 , n6694 );
and ( n8466 , n8465 , n6584 );
xor ( n8467 , n6584 , n6345 );
and ( n8468 , n8393 , n8394 );
xor ( n8469 , n8467 , n8468 );
and ( n8470 , n8469 , n6694 );
or ( n8471 , n8466 , n8470 );
and ( n8472 , n8471 , n5188 );
and ( n8473 , n4065 , n5282 );
or ( n8474 , n8472 , n8473 );
and ( n8475 , n8474 , n6710 );
and ( n8476 , n5529 , n5188 );
and ( n8477 , n4065 , n5282 );
or ( n8478 , n8476 , n8477 );
and ( n8479 , n8478 , n6717 );
and ( n8480 , n5529 , n6719 );
not ( n8481 , n5529 );
and ( n8482 , n8407 , n8408 );
xor ( n8483 , n8481 , n8482 );
and ( n8484 , n8483 , n5188 );
and ( n8485 , n4065 , n5282 );
or ( n8486 , n8484 , n8485 );
and ( n8487 , n8486 , n6724 );
or ( n8488 , n8426 , n8453 , n8464 , n8475 , n8479 , n8480 , n8487 );
and ( n8489 , n8425 , n8488 );
and ( n8490 , n4065 , n3260 );
or ( n8491 , n8489 , n8490 );
and ( n8492 , n8491 , n2422 );
and ( n8493 , n3860 , n2428 );
or ( n8494 , n8492 , n8493 );
buf ( n8495 , n8494 );
buf ( n8496 , n2424 );
buf ( n8497 , n2281 );
buf ( n8498 , n2280 );
not ( n8499 , n3260 );
and ( n8500 , n4055 , n3631 );
not ( n8501 , n7021 );
and ( n8502 , n8501 , n6939 );
xor ( n8503 , n6939 , n3770 );
and ( n8504 , n8429 , n8430 );
xor ( n8505 , n8503 , n8504 );
and ( n8506 , n8505 , n7021 );
or ( n8507 , n8502 , n8506 );
and ( n8508 , n8507 , n5289 );
and ( n8509 , n8507 , n5287 );
not ( n8510 , n3290 );
and ( n8511 , n8510 , n4884 );
not ( n8512 , n4999 );
and ( n8513 , n8512 , n4892 );
xor ( n8514 , n4892 , n4578 );
and ( n8515 , n8440 , n8441 );
xor ( n8516 , n8514 , n8515 );
and ( n8517 , n8516 , n4999 );
or ( n8518 , n8513 , n8517 );
and ( n8519 , n8518 , n3290 );
or ( n8520 , n8511 , n8519 );
and ( n8521 , n8520 , n5152 );
and ( n8522 , n4884 , n5154 );
or ( n8523 , n8508 , n8509 , n8521 , n8522 );
and ( n8524 , n8523 , n5188 );
and ( n8525 , n4055 , n5282 );
or ( n8526 , n8524 , n8525 );
and ( n8527 , n8526 , n5285 );
not ( n8528 , n6201 );
and ( n8529 , n8528 , n6103 );
xor ( n8530 , n6103 , n5852 );
and ( n8531 , n8456 , n8457 );
xor ( n8532 , n8530 , n8531 );
and ( n8533 , n8532 , n6201 );
or ( n8534 , n8529 , n8533 );
and ( n8535 , n8534 , n5188 );
and ( n8536 , n4055 , n5282 );
or ( n8537 , n8535 , n8536 );
and ( n8538 , n8537 , n6218 );
not ( n8539 , n6694 );
and ( n8540 , n8539 , n6596 );
xor ( n8541 , n6596 , n6345 );
and ( n8542 , n8467 , n8468 );
xor ( n8543 , n8541 , n8542 );
and ( n8544 , n8543 , n6694 );
or ( n8545 , n8540 , n8544 );
and ( n8546 , n8545 , n5188 );
and ( n8547 , n4055 , n5282 );
or ( n8548 , n8546 , n8547 );
and ( n8549 , n8548 , n6710 );
and ( n8550 , n5526 , n5188 );
and ( n8551 , n4055 , n5282 );
or ( n8552 , n8550 , n8551 );
and ( n8553 , n8552 , n6717 );
and ( n8554 , n5526 , n6719 );
not ( n8555 , n5526 );
and ( n8556 , n8481 , n8482 );
xor ( n8557 , n8555 , n8556 );
and ( n8558 , n8557 , n5188 );
and ( n8559 , n4055 , n5282 );
or ( n8560 , n8558 , n8559 );
and ( n8561 , n8560 , n6724 );
or ( n8562 , n8500 , n8527 , n8538 , n8549 , n8553 , n8554 , n8561 );
and ( n8563 , n8499 , n8562 );
and ( n8564 , n4055 , n3260 );
or ( n8565 , n8563 , n8564 );
and ( n8566 , n8565 , n2422 );
and ( n8567 , n3856 , n2428 );
or ( n8568 , n8566 , n8567 );
buf ( n8569 , n8568 );
buf ( n8570 , n2424 );
buf ( n8571 , n2281 );
buf ( n8572 , n2280 );
not ( n8573 , n3260 );
and ( n8574 , n4045 , n3631 );
not ( n8575 , n7021 );
and ( n8576 , n8575 , n6949 );
xor ( n8577 , n6949 , n3770 );
and ( n8578 , n8503 , n8504 );
xor ( n8579 , n8577 , n8578 );
and ( n8580 , n8579 , n7021 );
or ( n8581 , n8576 , n8580 );
and ( n8582 , n8581 , n5289 );
and ( n8583 , n8581 , n5287 );
not ( n8584 , n3290 );
and ( n8585 , n8584 , n4899 );
not ( n8586 , n4999 );
and ( n8587 , n8586 , n4907 );
xor ( n8588 , n4907 , n4578 );
and ( n8589 , n8514 , n8515 );
xor ( n8590 , n8588 , n8589 );
and ( n8591 , n8590 , n4999 );
or ( n8592 , n8587 , n8591 );
and ( n8593 , n8592 , n3290 );
or ( n8594 , n8585 , n8593 );
and ( n8595 , n8594 , n5152 );
and ( n8596 , n4899 , n5154 );
or ( n8597 , n8582 , n8583 , n8595 , n8596 );
and ( n8598 , n8597 , n5188 );
and ( n8599 , n4045 , n5282 );
or ( n8600 , n8598 , n8599 );
and ( n8601 , n8600 , n5285 );
not ( n8602 , n6201 );
and ( n8603 , n8602 , n6115 );
xor ( n8604 , n6115 , n5852 );
and ( n8605 , n8530 , n8531 );
xor ( n8606 , n8604 , n8605 );
and ( n8607 , n8606 , n6201 );
or ( n8608 , n8603 , n8607 );
and ( n8609 , n8608 , n5188 );
and ( n8610 , n4045 , n5282 );
or ( n8611 , n8609 , n8610 );
and ( n8612 , n8611 , n6218 );
not ( n8613 , n6694 );
and ( n8614 , n8613 , n6608 );
xor ( n8615 , n6608 , n6345 );
and ( n8616 , n8541 , n8542 );
xor ( n8617 , n8615 , n8616 );
and ( n8618 , n8617 , n6694 );
or ( n8619 , n8614 , n8618 );
and ( n8620 , n8619 , n5188 );
and ( n8621 , n4045 , n5282 );
or ( n8622 , n8620 , n8621 );
and ( n8623 , n8622 , n6710 );
and ( n8624 , n5523 , n5188 );
and ( n8625 , n4045 , n5282 );
or ( n8626 , n8624 , n8625 );
and ( n8627 , n8626 , n6717 );
and ( n8628 , n5523 , n6719 );
not ( n8629 , n5523 );
and ( n8630 , n8555 , n8556 );
xor ( n8631 , n8629 , n8630 );
and ( n8632 , n8631 , n5188 );
and ( n8633 , n4045 , n5282 );
or ( n8634 , n8632 , n8633 );
and ( n8635 , n8634 , n6724 );
or ( n8636 , n8574 , n8601 , n8612 , n8623 , n8627 , n8628 , n8635 );
and ( n8637 , n8573 , n8636 );
and ( n8638 , n4045 , n3260 );
or ( n8639 , n8637 , n8638 );
and ( n8640 , n8639 , n2422 );
and ( n8641 , n3851 , n2428 );
or ( n8642 , n8640 , n8641 );
buf ( n8643 , n8642 );
buf ( n8644 , n2424 );
buf ( n8645 , n2281 );
buf ( n8646 , n2280 );
not ( n8647 , n3260 );
and ( n8648 , n4035 , n3631 );
not ( n8649 , n7021 );
and ( n8650 , n8649 , n6959 );
xor ( n8651 , n6959 , n3770 );
and ( n8652 , n8577 , n8578 );
xor ( n8653 , n8651 , n8652 );
and ( n8654 , n8653 , n7021 );
or ( n8655 , n8650 , n8654 );
and ( n8656 , n8655 , n5289 );
and ( n8657 , n8655 , n5287 );
not ( n8658 , n3290 );
and ( n8659 , n8658 , n4914 );
not ( n8660 , n4999 );
and ( n8661 , n8660 , n4922 );
xor ( n8662 , n4922 , n4578 );
and ( n8663 , n8588 , n8589 );
xor ( n8664 , n8662 , n8663 );
and ( n8665 , n8664 , n4999 );
or ( n8666 , n8661 , n8665 );
and ( n8667 , n8666 , n3290 );
or ( n8668 , n8659 , n8667 );
and ( n8669 , n8668 , n5152 );
and ( n8670 , n4914 , n5154 );
or ( n8671 , n8656 , n8657 , n8669 , n8670 );
and ( n8672 , n8671 , n5188 );
and ( n8673 , n4035 , n5282 );
or ( n8674 , n8672 , n8673 );
and ( n8675 , n8674 , n5285 );
not ( n8676 , n6201 );
and ( n8677 , n8676 , n6127 );
xor ( n8678 , n6127 , n5852 );
and ( n8679 , n8604 , n8605 );
xor ( n8680 , n8678 , n8679 );
and ( n8681 , n8680 , n6201 );
or ( n8682 , n8677 , n8681 );
and ( n8683 , n8682 , n5188 );
and ( n8684 , n4035 , n5282 );
or ( n8685 , n8683 , n8684 );
and ( n8686 , n8685 , n6218 );
not ( n8687 , n6694 );
and ( n8688 , n8687 , n6620 );
xor ( n8689 , n6620 , n6345 );
and ( n8690 , n8615 , n8616 );
xor ( n8691 , n8689 , n8690 );
and ( n8692 , n8691 , n6694 );
or ( n8693 , n8688 , n8692 );
and ( n8694 , n8693 , n5188 );
and ( n8695 , n4035 , n5282 );
or ( n8696 , n8694 , n8695 );
and ( n8697 , n8696 , n6710 );
and ( n8698 , n5520 , n5188 );
and ( n8699 , n4035 , n5282 );
or ( n8700 , n8698 , n8699 );
and ( n8701 , n8700 , n6717 );
and ( n8702 , n5520 , n6719 );
not ( n8703 , n5520 );
and ( n8704 , n8629 , n8630 );
xor ( n8705 , n8703 , n8704 );
and ( n8706 , n8705 , n5188 );
and ( n8707 , n4035 , n5282 );
or ( n8708 , n8706 , n8707 );
and ( n8709 , n8708 , n6724 );
or ( n8710 , n8648 , n8675 , n8686 , n8697 , n8701 , n8702 , n8709 );
and ( n8711 , n8647 , n8710 );
and ( n8712 , n4035 , n3260 );
or ( n8713 , n8711 , n8712 );
and ( n8714 , n8713 , n2422 );
and ( n8715 , n3846 , n2428 );
or ( n8716 , n8714 , n8715 );
buf ( n8717 , n8716 );
buf ( n8718 , n2424 );
buf ( n8719 , n2281 );
buf ( n8720 , n2280 );
not ( n8721 , n3260 );
and ( n8722 , n4025 , n3631 );
not ( n8723 , n7021 );
and ( n8724 , n8723 , n6969 );
xor ( n8725 , n6969 , n3770 );
and ( n8726 , n8651 , n8652 );
xor ( n8727 , n8725 , n8726 );
and ( n8728 , n8727 , n7021 );
or ( n8729 , n8724 , n8728 );
and ( n8730 , n8729 , n5289 );
and ( n8731 , n8729 , n5287 );
not ( n8732 , n3290 );
and ( n8733 , n8732 , n4929 );
not ( n8734 , n4999 );
and ( n8735 , n8734 , n4937 );
xor ( n8736 , n4937 , n4578 );
and ( n8737 , n8662 , n8663 );
xor ( n8738 , n8736 , n8737 );
and ( n8739 , n8738 , n4999 );
or ( n8740 , n8735 , n8739 );
and ( n8741 , n8740 , n3290 );
or ( n8742 , n8733 , n8741 );
and ( n8743 , n8742 , n5152 );
and ( n8744 , n4929 , n5154 );
or ( n8745 , n8730 , n8731 , n8743 , n8744 );
and ( n8746 , n8745 , n5188 );
and ( n8747 , n4025 , n5282 );
or ( n8748 , n8746 , n8747 );
and ( n8749 , n8748 , n5285 );
not ( n8750 , n6201 );
and ( n8751 , n8750 , n6139 );
xor ( n8752 , n6139 , n5852 );
and ( n8753 , n8678 , n8679 );
xor ( n8754 , n8752 , n8753 );
and ( n8755 , n8754 , n6201 );
or ( n8756 , n8751 , n8755 );
and ( n8757 , n8756 , n5188 );
and ( n8758 , n4025 , n5282 );
or ( n8759 , n8757 , n8758 );
and ( n8760 , n8759 , n6218 );
not ( n8761 , n6694 );
and ( n8762 , n8761 , n6632 );
xor ( n8763 , n6632 , n6345 );
and ( n8764 , n8689 , n8690 );
xor ( n8765 , n8763 , n8764 );
and ( n8766 , n8765 , n6694 );
or ( n8767 , n8762 , n8766 );
and ( n8768 , n8767 , n5188 );
and ( n8769 , n4025 , n5282 );
or ( n8770 , n8768 , n8769 );
and ( n8771 , n8770 , n6710 );
and ( n8772 , n5517 , n5188 );
and ( n8773 , n4025 , n5282 );
or ( n8774 , n8772 , n8773 );
and ( n8775 , n8774 , n6717 );
and ( n8776 , n5517 , n6719 );
not ( n8777 , n5517 );
and ( n8778 , n8703 , n8704 );
xor ( n8779 , n8777 , n8778 );
and ( n8780 , n8779 , n5188 );
and ( n8781 , n4025 , n5282 );
or ( n8782 , n8780 , n8781 );
and ( n8783 , n8782 , n6724 );
or ( n8784 , n8722 , n8749 , n8760 , n8771 , n8775 , n8776 , n8783 );
and ( n8785 , n8721 , n8784 );
and ( n8786 , n4025 , n3260 );
or ( n8787 , n8785 , n8786 );
and ( n8788 , n8787 , n2422 );
and ( n8789 , n3841 , n2428 );
or ( n8790 , n8788 , n8789 );
buf ( n8791 , n8790 );
buf ( n8792 , n2424 );
buf ( n8793 , n2281 );
buf ( n8794 , n2280 );
not ( n8795 , n3260 );
and ( n8796 , n4015 , n3631 );
not ( n8797 , n7021 );
and ( n8798 , n8797 , n6979 );
xor ( n8799 , n6979 , n3770 );
and ( n8800 , n8725 , n8726 );
xor ( n8801 , n8799 , n8800 );
and ( n8802 , n8801 , n7021 );
or ( n8803 , n8798 , n8802 );
and ( n8804 , n8803 , n5289 );
and ( n8805 , n8803 , n5287 );
not ( n8806 , n3290 );
and ( n8807 , n8806 , n4944 );
not ( n8808 , n4999 );
and ( n8809 , n8808 , n4952 );
xor ( n8810 , n4952 , n4578 );
and ( n8811 , n8736 , n8737 );
xor ( n8812 , n8810 , n8811 );
and ( n8813 , n8812 , n4999 );
or ( n8814 , n8809 , n8813 );
and ( n8815 , n8814 , n3290 );
or ( n8816 , n8807 , n8815 );
and ( n8817 , n8816 , n5152 );
and ( n8818 , n4944 , n5154 );
or ( n8819 , n8804 , n8805 , n8817 , n8818 );
and ( n8820 , n8819 , n5188 );
and ( n8821 , n4015 , n5282 );
or ( n8822 , n8820 , n8821 );
and ( n8823 , n8822 , n5285 );
not ( n8824 , n6201 );
and ( n8825 , n8824 , n6151 );
xor ( n8826 , n6151 , n5852 );
and ( n8827 , n8752 , n8753 );
xor ( n8828 , n8826 , n8827 );
and ( n8829 , n8828 , n6201 );
or ( n8830 , n8825 , n8829 );
and ( n8831 , n8830 , n5188 );
and ( n8832 , n4015 , n5282 );
or ( n8833 , n8831 , n8832 );
and ( n8834 , n8833 , n6218 );
not ( n8835 , n6694 );
and ( n8836 , n8835 , n6644 );
xor ( n8837 , n6644 , n6345 );
and ( n8838 , n8763 , n8764 );
xor ( n8839 , n8837 , n8838 );
and ( n8840 , n8839 , n6694 );
or ( n8841 , n8836 , n8840 );
and ( n8842 , n8841 , n5188 );
and ( n8843 , n4015 , n5282 );
or ( n8844 , n8842 , n8843 );
and ( n8845 , n8844 , n6710 );
and ( n8846 , n5514 , n5188 );
and ( n8847 , n4015 , n5282 );
or ( n8848 , n8846 , n8847 );
and ( n8849 , n8848 , n6717 );
and ( n8850 , n5514 , n6719 );
not ( n8851 , n5514 );
and ( n8852 , n8777 , n8778 );
xor ( n8853 , n8851 , n8852 );
and ( n8854 , n8853 , n5188 );
and ( n8855 , n4015 , n5282 );
or ( n8856 , n8854 , n8855 );
and ( n8857 , n8856 , n6724 );
or ( n8858 , n8796 , n8823 , n8834 , n8845 , n8849 , n8850 , n8857 );
and ( n8859 , n8795 , n8858 );
and ( n8860 , n4015 , n3260 );
or ( n8861 , n8859 , n8860 );
and ( n8862 , n8861 , n2422 );
and ( n8863 , n3836 , n2428 );
or ( n8864 , n8862 , n8863 );
buf ( n8865 , n8864 );
buf ( n8866 , n2424 );
buf ( n8867 , n2281 );
buf ( n8868 , n2280 );
not ( n8869 , n3260 );
and ( n8870 , n4005 , n3631 );
not ( n8871 , n7021 );
and ( n8872 , n8871 , n6989 );
xor ( n8873 , n6989 , n3770 );
and ( n8874 , n8799 , n8800 );
xor ( n8875 , n8873 , n8874 );
and ( n8876 , n8875 , n7021 );
or ( n8877 , n8872 , n8876 );
and ( n8878 , n8877 , n5289 );
and ( n8879 , n8877 , n5287 );
not ( n8880 , n3290 );
and ( n8881 , n8880 , n4959 );
not ( n8882 , n4999 );
and ( n8883 , n8882 , n4967 );
xor ( n8884 , n4967 , n4578 );
and ( n8885 , n8810 , n8811 );
xor ( n8886 , n8884 , n8885 );
and ( n8887 , n8886 , n4999 );
or ( n8888 , n8883 , n8887 );
and ( n8889 , n8888 , n3290 );
or ( n8890 , n8881 , n8889 );
and ( n8891 , n8890 , n5152 );
and ( n8892 , n4959 , n5154 );
or ( n8893 , n8878 , n8879 , n8891 , n8892 );
and ( n8894 , n8893 , n5188 );
and ( n8895 , n4005 , n5282 );
or ( n8896 , n8894 , n8895 );
and ( n8897 , n8896 , n5285 );
not ( n8898 , n6201 );
and ( n8899 , n8898 , n6163 );
xor ( n8900 , n6163 , n5852 );
and ( n8901 , n8826 , n8827 );
xor ( n8902 , n8900 , n8901 );
and ( n8903 , n8902 , n6201 );
or ( n8904 , n8899 , n8903 );
and ( n8905 , n8904 , n5188 );
and ( n8906 , n4005 , n5282 );
or ( n8907 , n8905 , n8906 );
and ( n8908 , n8907 , n6218 );
not ( n8909 , n6694 );
and ( n8910 , n8909 , n6656 );
xor ( n8911 , n6656 , n6345 );
and ( n8912 , n8837 , n8838 );
xor ( n8913 , n8911 , n8912 );
and ( n8914 , n8913 , n6694 );
or ( n8915 , n8910 , n8914 );
and ( n8916 , n8915 , n5188 );
and ( n8917 , n4005 , n5282 );
or ( n8918 , n8916 , n8917 );
and ( n8919 , n8918 , n6710 );
and ( n8920 , n5511 , n5188 );
and ( n8921 , n4005 , n5282 );
or ( n8922 , n8920 , n8921 );
and ( n8923 , n8922 , n6717 );
and ( n8924 , n5511 , n6719 );
not ( n8925 , n5511 );
and ( n8926 , n8851 , n8852 );
xor ( n8927 , n8925 , n8926 );
and ( n8928 , n8927 , n5188 );
and ( n8929 , n4005 , n5282 );
or ( n8930 , n8928 , n8929 );
and ( n8931 , n8930 , n6724 );
or ( n8932 , n8870 , n8897 , n8908 , n8919 , n8923 , n8924 , n8931 );
and ( n8933 , n8869 , n8932 );
and ( n8934 , n4005 , n3260 );
or ( n8935 , n8933 , n8934 );
and ( n8936 , n8935 , n2422 );
and ( n8937 , n3831 , n2428 );
or ( n8938 , n8936 , n8937 );
buf ( n8939 , n8938 );
buf ( n8940 , n2424 );
buf ( n8941 , n2281 );
buf ( n8942 , n2280 );
not ( n8943 , n3260 );
and ( n8944 , n3995 , n3631 );
not ( n8945 , n7021 );
and ( n8946 , n8945 , n6999 );
xor ( n8947 , n6999 , n3770 );
and ( n8948 , n8873 , n8874 );
xor ( n8949 , n8947 , n8948 );
and ( n8950 , n8949 , n7021 );
or ( n8951 , n8946 , n8950 );
and ( n8952 , n8951 , n5289 );
and ( n8953 , n8951 , n5287 );
not ( n8954 , n3290 );
and ( n8955 , n8954 , n4974 );
not ( n8956 , n4999 );
and ( n8957 , n8956 , n4982 );
xor ( n8958 , n4982 , n4578 );
and ( n8959 , n8884 , n8885 );
xor ( n8960 , n8958 , n8959 );
and ( n8961 , n8960 , n4999 );
or ( n8962 , n8957 , n8961 );
and ( n8963 , n8962 , n3290 );
or ( n8964 , n8955 , n8963 );
and ( n8965 , n8964 , n5152 );
and ( n8966 , n4974 , n5154 );
or ( n8967 , n8952 , n8953 , n8965 , n8966 );
and ( n8968 , n8967 , n5188 );
and ( n8969 , n3995 , n5282 );
or ( n8970 , n8968 , n8969 );
and ( n8971 , n8970 , n5285 );
not ( n8972 , n6201 );
and ( n8973 , n8972 , n6175 );
xor ( n8974 , n6175 , n5852 );
and ( n8975 , n8900 , n8901 );
xor ( n8976 , n8974 , n8975 );
and ( n8977 , n8976 , n6201 );
or ( n8978 , n8973 , n8977 );
and ( n8979 , n8978 , n5188 );
and ( n8980 , n3995 , n5282 );
or ( n8981 , n8979 , n8980 );
and ( n8982 , n8981 , n6218 );
not ( n8983 , n6694 );
and ( n8984 , n8983 , n6668 );
xor ( n8985 , n6668 , n6345 );
and ( n8986 , n8911 , n8912 );
xor ( n8987 , n8985 , n8986 );
and ( n8988 , n8987 , n6694 );
or ( n8989 , n8984 , n8988 );
and ( n8990 , n8989 , n5188 );
and ( n8991 , n3995 , n5282 );
or ( n8992 , n8990 , n8991 );
and ( n8993 , n8992 , n6710 );
and ( n8994 , n5508 , n5188 );
and ( n8995 , n3995 , n5282 );
or ( n8996 , n8994 , n8995 );
and ( n8997 , n8996 , n6717 );
and ( n8998 , n5508 , n6719 );
not ( n8999 , n5508 );
and ( n9000 , n8925 , n8926 );
xor ( n9001 , n8999 , n9000 );
and ( n9002 , n9001 , n5188 );
and ( n9003 , n3995 , n5282 );
or ( n9004 , n9002 , n9003 );
and ( n9005 , n9004 , n6724 );
or ( n9006 , n8944 , n8971 , n8982 , n8993 , n8997 , n8998 , n9005 );
and ( n9007 , n8943 , n9006 );
and ( n9008 , n3995 , n3260 );
or ( n9009 , n9007 , n9008 );
and ( n9010 , n9009 , n2422 );
and ( n9011 , n3826 , n2428 );
or ( n9012 , n9010 , n9011 );
buf ( n9013 , n9012 );
buf ( n9014 , n2424 );
buf ( n9015 , n2281 );
buf ( n9016 , n2280 );
not ( n9017 , n3260 );
and ( n9018 , n3985 , n3631 );
not ( n9019 , n7021 );
and ( n9020 , n9019 , n7009 );
xor ( n9021 , n7009 , n3770 );
and ( n9022 , n8947 , n8948 );
xor ( n9023 , n9021 , n9022 );
and ( n9024 , n9023 , n7021 );
or ( n9025 , n9020 , n9024 );
and ( n9026 , n9025 , n5289 );
and ( n9027 , n9025 , n5287 );
not ( n9028 , n3290 );
and ( n9029 , n9028 , n4989 );
not ( n9030 , n4999 );
and ( n9031 , n9030 , n4997 );
xor ( n9032 , n4997 , n4578 );
and ( n9033 , n8958 , n8959 );
xor ( n9034 , n9032 , n9033 );
and ( n9035 , n9034 , n4999 );
or ( n9036 , n9031 , n9035 );
and ( n9037 , n9036 , n3290 );
or ( n9038 , n9029 , n9037 );
and ( n9039 , n9038 , n5152 );
and ( n9040 , n4989 , n5154 );
or ( n9041 , n9026 , n9027 , n9039 , n9040 );
and ( n9042 , n9041 , n5188 );
and ( n9043 , n3985 , n5282 );
or ( n9044 , n9042 , n9043 );
and ( n9045 , n9044 , n5285 );
not ( n9046 , n6201 );
and ( n9047 , n9046 , n6187 );
xor ( n9048 , n6187 , n5852 );
and ( n9049 , n8974 , n8975 );
xor ( n9050 , n9048 , n9049 );
and ( n9051 , n9050 , n6201 );
or ( n9052 , n9047 , n9051 );
and ( n9053 , n9052 , n5188 );
and ( n9054 , n3985 , n5282 );
or ( n9055 , n9053 , n9054 );
and ( n9056 , n9055 , n6218 );
not ( n9057 , n6694 );
and ( n9058 , n9057 , n6680 );
xor ( n9059 , n6680 , n6345 );
and ( n9060 , n8985 , n8986 );
xor ( n9061 , n9059 , n9060 );
and ( n9062 , n9061 , n6694 );
or ( n9063 , n9058 , n9062 );
and ( n9064 , n9063 , n5188 );
and ( n9065 , n3985 , n5282 );
or ( n9066 , n9064 , n9065 );
and ( n9067 , n9066 , n6710 );
and ( n9068 , n5505 , n5188 );
and ( n9069 , n3985 , n5282 );
or ( n9070 , n9068 , n9069 );
and ( n9071 , n9070 , n6717 );
and ( n9072 , n5505 , n6719 );
not ( n9073 , n5505 );
and ( n9074 , n8999 , n9000 );
xor ( n9075 , n9073 , n9074 );
and ( n9076 , n9075 , n5188 );
and ( n9077 , n3985 , n5282 );
or ( n9078 , n9076 , n9077 );
and ( n9079 , n9078 , n6724 );
or ( n9080 , n9018 , n9045 , n9056 , n9067 , n9071 , n9072 , n9079 );
and ( n9081 , n9017 , n9080 );
and ( n9082 , n3985 , n3260 );
or ( n9083 , n9081 , n9082 );
and ( n9084 , n9083 , n2422 );
and ( n9085 , n3821 , n2428 );
or ( n9086 , n9084 , n9085 );
buf ( n9087 , n9086 );
buf ( n9088 , n2424 );
buf ( n9089 , n2281 );
buf ( n9090 , n2280 );
not ( n9091 , n3260 );
and ( n9092 , n5156 , n5219 );
or ( n9093 , n5249 , n5280 );
or ( n9094 , n9093 , n5188 );
buf ( n9095 , n9094 );
and ( n9096 , n3791 , n9095 );
or ( n9097 , n9092 , n9096 );
and ( n9098 , n9097 , n5285 );
and ( n9099 , n6207 , n5219 );
and ( n9100 , n3791 , n9095 );
or ( n9101 , n9099 , n9100 );
and ( n9102 , n9101 , n6218 );
and ( n9103 , n6700 , n5219 );
and ( n9104 , n3791 , n9095 );
or ( n9105 , n9103 , n9104 );
and ( n9106 , n9105 , n6710 );
and ( n9107 , n5492 , n5219 );
and ( n9108 , n3791 , n9095 );
or ( n9109 , n9107 , n9108 );
and ( n9110 , n9109 , n6717 );
and ( n9111 , n5492 , n5219 );
and ( n9112 , n3791 , n9095 );
or ( n9113 , n9111 , n9112 );
and ( n9114 , n9113 , n6724 );
or ( n9115 , n6719 , n3631 );
and ( n9116 , n3791 , n9115 );
or ( n9117 , n9098 , n9102 , n9106 , n9110 , n9114 , n9116 );
and ( n9118 , n9091 , n9117 );
and ( n9119 , n3791 , n3260 );
or ( n9120 , n9118 , n9119 );
and ( n9121 , n9120 , n2422 );
and ( n9122 , n3791 , n2428 );
or ( n9123 , n9121 , n9122 );
buf ( n9124 , n9123 );
buf ( n9125 , n2424 );
buf ( n9126 , n2281 );
buf ( n9127 , n2280 );
not ( n9128 , n3260 );
and ( n9129 , n7043 , n5219 );
and ( n9130 , n3781 , n9095 );
or ( n9131 , n9129 , n9130 );
and ( n9132 , n9131 , n5285 );
and ( n9133 , n7054 , n5219 );
and ( n9134 , n3781 , n9095 );
or ( n9135 , n9133 , n9134 );
and ( n9136 , n9135 , n6218 );
and ( n9137 , n7065 , n5219 );
and ( n9138 , n3781 , n9095 );
or ( n9139 , n9137 , n9138 );
and ( n9140 , n9139 , n6710 );
and ( n9141 , n5757 , n5219 );
and ( n9142 , n3781 , n9095 );
or ( n9143 , n9141 , n9142 );
and ( n9144 , n9143 , n6717 );
and ( n9145 , n7077 , n5219 );
and ( n9146 , n3781 , n9095 );
or ( n9147 , n9145 , n9146 );
and ( n9148 , n9147 , n6724 );
and ( n9149 , n3781 , n9115 );
or ( n9150 , n9132 , n9136 , n9140 , n9144 , n9148 , n9149 );
and ( n9151 , n9128 , n9150 );
and ( n9152 , n3781 , n3260 );
or ( n9153 , n9151 , n9152 );
and ( n9154 , n9153 , n2422 );
and ( n9155 , n3781 , n2428 );
or ( n9156 , n9154 , n9155 );
buf ( n9157 , n9156 );
buf ( n9158 , n2424 );
buf ( n9159 , n2281 );
buf ( n9160 , n2280 );
not ( n9161 , n3260 );
and ( n9162 , n7117 , n5219 );
and ( n9163 , n4253 , n9095 );
or ( n9164 , n9162 , n9163 );
and ( n9165 , n9164 , n5285 );
and ( n9166 , n7128 , n5219 );
and ( n9167 , n4253 , n9095 );
or ( n9168 , n9166 , n9167 );
and ( n9169 , n9168 , n6218 );
and ( n9170 , n7139 , n5219 );
and ( n9171 , n4253 , n9095 );
or ( n9172 , n9170 , n9171 );
and ( n9173 , n9172 , n6710 );
and ( n9174 , n5747 , n5219 );
and ( n9175 , n4253 , n9095 );
or ( n9176 , n9174 , n9175 );
and ( n9177 , n9176 , n6717 );
and ( n9178 , n7151 , n5219 );
and ( n9179 , n4253 , n9095 );
or ( n9180 , n9178 , n9179 );
and ( n9181 , n9180 , n6724 );
and ( n9182 , n4253 , n9115 );
or ( n9183 , n9165 , n9169 , n9173 , n9177 , n9181 , n9182 );
and ( n9184 , n9161 , n9183 );
and ( n9185 , n4253 , n3260 );
or ( n9186 , n9184 , n9185 );
and ( n9187 , n9186 , n2422 );
and ( n9188 , n4253 , n2428 );
or ( n9189 , n9187 , n9188 );
buf ( n9190 , n9189 );
buf ( n9191 , n2424 );
buf ( n9192 , n2281 );
buf ( n9193 , n2280 );
not ( n9194 , n3260 );
and ( n9195 , n7191 , n5219 );
and ( n9196 , n4239 , n9095 );
or ( n9197 , n9195 , n9196 );
and ( n9198 , n9197 , n5285 );
and ( n9199 , n7202 , n5219 );
and ( n9200 , n4239 , n9095 );
or ( n9201 , n9199 , n9200 );
and ( n9202 , n9201 , n6218 );
and ( n9203 , n7213 , n5219 );
and ( n9204 , n4239 , n9095 );
or ( n9205 , n9203 , n9204 );
and ( n9206 , n9205 , n6710 );
and ( n9207 , n5737 , n5219 );
and ( n9208 , n4239 , n9095 );
or ( n9209 , n9207 , n9208 );
and ( n9210 , n9209 , n6717 );
and ( n9211 , n7225 , n5219 );
and ( n9212 , n4239 , n9095 );
or ( n9213 , n9211 , n9212 );
and ( n9214 , n9213 , n6724 );
and ( n9215 , n4239 , n9115 );
or ( n9216 , n9198 , n9202 , n9206 , n9210 , n9214 , n9215 );
and ( n9217 , n9194 , n9216 );
and ( n9218 , n4239 , n3260 );
or ( n9219 , n9217 , n9218 );
and ( n9220 , n9219 , n2422 );
and ( n9221 , n4239 , n2428 );
or ( n9222 , n9220 , n9221 );
buf ( n9223 , n9222 );
buf ( n9224 , n2424 );
buf ( n9225 , n2281 );
buf ( n9226 , n2280 );
not ( n9227 , n3260 );
and ( n9228 , n7265 , n5219 );
and ( n9229 , n4229 , n9095 );
or ( n9230 , n9228 , n9229 );
and ( n9231 , n9230 , n5285 );
and ( n9232 , n7276 , n5219 );
and ( n9233 , n4229 , n9095 );
or ( n9234 , n9232 , n9233 );
and ( n9235 , n9234 , n6218 );
and ( n9236 , n7287 , n5219 );
and ( n9237 , n4229 , n9095 );
or ( n9238 , n9236 , n9237 );
and ( n9239 , n9238 , n6710 );
and ( n9240 , n5727 , n5219 );
and ( n9241 , n4229 , n9095 );
or ( n9242 , n9240 , n9241 );
and ( n9243 , n9242 , n6717 );
and ( n9244 , n7299 , n5219 );
and ( n9245 , n4229 , n9095 );
or ( n9246 , n9244 , n9245 );
and ( n9247 , n9246 , n6724 );
and ( n9248 , n4229 , n9115 );
or ( n9249 , n9231 , n9235 , n9239 , n9243 , n9247 , n9248 );
and ( n9250 , n9227 , n9249 );
and ( n9251 , n4229 , n3260 );
or ( n9252 , n9250 , n9251 );
and ( n9253 , n9252 , n2422 );
and ( n9254 , n4229 , n2428 );
or ( n9255 , n9253 , n9254 );
buf ( n9256 , n9255 );
buf ( n9257 , n2424 );
buf ( n9258 , n2281 );
buf ( n9259 , n2280 );
not ( n9260 , n3260 );
and ( n9261 , n7339 , n5219 );
and ( n9262 , n4219 , n9095 );
or ( n9263 , n9261 , n9262 );
and ( n9264 , n9263 , n5285 );
and ( n9265 , n7350 , n5219 );
and ( n9266 , n4219 , n9095 );
or ( n9267 , n9265 , n9266 );
and ( n9268 , n9267 , n6218 );
and ( n9269 , n7361 , n5219 );
and ( n9270 , n4219 , n9095 );
or ( n9271 , n9269 , n9270 );
and ( n9272 , n9271 , n6710 );
and ( n9273 , n5717 , n5219 );
and ( n9274 , n4219 , n9095 );
or ( n9275 , n9273 , n9274 );
and ( n9276 , n9275 , n6717 );
and ( n9277 , n7373 , n5219 );
and ( n9278 , n4219 , n9095 );
or ( n9279 , n9277 , n9278 );
and ( n9280 , n9279 , n6724 );
and ( n9281 , n4219 , n9115 );
or ( n9282 , n9264 , n9268 , n9272 , n9276 , n9280 , n9281 );
and ( n9283 , n9260 , n9282 );
and ( n9284 , n4219 , n3260 );
or ( n9285 , n9283 , n9284 );
and ( n9286 , n9285 , n2422 );
and ( n9287 , n4219 , n2428 );
or ( n9288 , n9286 , n9287 );
buf ( n9289 , n9288 );
buf ( n9290 , n2424 );
buf ( n9291 , n2281 );
buf ( n9292 , n2280 );
not ( n9293 , n3260 );
and ( n9294 , n7413 , n5219 );
and ( n9295 , n4209 , n9095 );
or ( n9296 , n9294 , n9295 );
and ( n9297 , n9296 , n5285 );
and ( n9298 , n7424 , n5219 );
and ( n9299 , n4209 , n9095 );
or ( n9300 , n9298 , n9299 );
and ( n9301 , n9300 , n6218 );
and ( n9302 , n7435 , n5219 );
and ( n9303 , n4209 , n9095 );
or ( n9304 , n9302 , n9303 );
and ( n9305 , n9304 , n6710 );
and ( n9306 , n5707 , n5219 );
and ( n9307 , n4209 , n9095 );
or ( n9308 , n9306 , n9307 );
and ( n9309 , n9308 , n6717 );
and ( n9310 , n7447 , n5219 );
and ( n9311 , n4209 , n9095 );
or ( n9312 , n9310 , n9311 );
and ( n9313 , n9312 , n6724 );
and ( n9314 , n4209 , n9115 );
or ( n9315 , n9297 , n9301 , n9305 , n9309 , n9313 , n9314 );
and ( n9316 , n9293 , n9315 );
and ( n9317 , n4209 , n3260 );
or ( n9318 , n9316 , n9317 );
and ( n9319 , n9318 , n2422 );
and ( n9320 , n4209 , n2428 );
or ( n9321 , n9319 , n9320 );
buf ( n9322 , n9321 );
buf ( n9323 , n2424 );
buf ( n9324 , n2281 );
buf ( n9325 , n2280 );
not ( n9326 , n3260 );
and ( n9327 , n7487 , n5219 );
and ( n9328 , n4199 , n9095 );
or ( n9329 , n9327 , n9328 );
and ( n9330 , n9329 , n5285 );
and ( n9331 , n7498 , n5219 );
and ( n9332 , n4199 , n9095 );
or ( n9333 , n9331 , n9332 );
and ( n9334 , n9333 , n6218 );
and ( n9335 , n7509 , n5219 );
and ( n9336 , n4199 , n9095 );
or ( n9337 , n9335 , n9336 );
and ( n9338 , n9337 , n6710 );
and ( n9339 , n5697 , n5219 );
and ( n9340 , n4199 , n9095 );
or ( n9341 , n9339 , n9340 );
and ( n9342 , n9341 , n6717 );
and ( n9343 , n7521 , n5219 );
and ( n9344 , n4199 , n9095 );
or ( n9345 , n9343 , n9344 );
and ( n9346 , n9345 , n6724 );
and ( n9347 , n4199 , n9115 );
or ( n9348 , n9330 , n9334 , n9338 , n9342 , n9346 , n9347 );
and ( n9349 , n9326 , n9348 );
and ( n9350 , n4199 , n3260 );
or ( n9351 , n9349 , n9350 );
and ( n9352 , n9351 , n2422 );
and ( n9353 , n4199 , n2428 );
or ( n9354 , n9352 , n9353 );
buf ( n9355 , n9354 );
buf ( n9356 , n2424 );
buf ( n9357 , n2281 );
buf ( n9358 , n2280 );
not ( n9359 , n3260 );
and ( n9360 , n7561 , n5219 );
and ( n9361 , n4189 , n9095 );
or ( n9362 , n9360 , n9361 );
and ( n9363 , n9362 , n5285 );
and ( n9364 , n7572 , n5219 );
and ( n9365 , n4189 , n9095 );
or ( n9366 , n9364 , n9365 );
and ( n9367 , n9366 , n6218 );
and ( n9368 , n7583 , n5219 );
and ( n9369 , n4189 , n9095 );
or ( n9370 , n9368 , n9369 );
and ( n9371 , n9370 , n6710 );
and ( n9372 , n5687 , n5219 );
and ( n9373 , n4189 , n9095 );
or ( n9374 , n9372 , n9373 );
and ( n9375 , n9374 , n6717 );
and ( n9376 , n7595 , n5219 );
and ( n9377 , n4189 , n9095 );
or ( n9378 , n9376 , n9377 );
and ( n9379 , n9378 , n6724 );
and ( n9380 , n4189 , n9115 );
or ( n9381 , n9363 , n9367 , n9371 , n9375 , n9379 , n9380 );
and ( n9382 , n9359 , n9381 );
and ( n9383 , n4189 , n3260 );
or ( n9384 , n9382 , n9383 );
and ( n9385 , n9384 , n2422 );
and ( n9386 , n4189 , n2428 );
or ( n9387 , n9385 , n9386 );
buf ( n9388 , n9387 );
buf ( n9389 , n2424 );
buf ( n9390 , n2281 );
buf ( n9391 , n2280 );
not ( n9392 , n3260 );
and ( n9393 , n7635 , n5219 );
and ( n9394 , n4179 , n9095 );
or ( n9395 , n9393 , n9394 );
and ( n9396 , n9395 , n5285 );
and ( n9397 , n7646 , n5219 );
and ( n9398 , n4179 , n9095 );
or ( n9399 , n9397 , n9398 );
and ( n9400 , n9399 , n6218 );
and ( n9401 , n7657 , n5219 );
and ( n9402 , n4179 , n9095 );
or ( n9403 , n9401 , n9402 );
and ( n9404 , n9403 , n6710 );
and ( n9405 , n5677 , n5219 );
and ( n9406 , n4179 , n9095 );
or ( n9407 , n9405 , n9406 );
and ( n9408 , n9407 , n6717 );
and ( n9409 , n7669 , n5219 );
and ( n9410 , n4179 , n9095 );
or ( n9411 , n9409 , n9410 );
and ( n9412 , n9411 , n6724 );
and ( n9413 , n4179 , n9115 );
or ( n9414 , n9396 , n9400 , n9404 , n9408 , n9412 , n9413 );
and ( n9415 , n9392 , n9414 );
and ( n9416 , n4179 , n3260 );
or ( n9417 , n9415 , n9416 );
and ( n9418 , n9417 , n2422 );
and ( n9419 , n4179 , n2428 );
or ( n9420 , n9418 , n9419 );
buf ( n9421 , n9420 );
buf ( n9422 , n2424 );
buf ( n9423 , n2281 );
buf ( n9424 , n2280 );
not ( n9425 , n3260 );
and ( n9426 , n7709 , n5219 );
and ( n9427 , n4169 , n9095 );
or ( n9428 , n9426 , n9427 );
and ( n9429 , n9428 , n5285 );
and ( n9430 , n7720 , n5219 );
and ( n9431 , n4169 , n9095 );
or ( n9432 , n9430 , n9431 );
and ( n9433 , n9432 , n6218 );
and ( n9434 , n7731 , n5219 );
and ( n9435 , n4169 , n9095 );
or ( n9436 , n9434 , n9435 );
and ( n9437 , n9436 , n6710 );
and ( n9438 , n5667 , n5219 );
and ( n9439 , n4169 , n9095 );
or ( n9440 , n9438 , n9439 );
and ( n9441 , n9440 , n6717 );
and ( n9442 , n7743 , n5219 );
and ( n9443 , n4169 , n9095 );
or ( n9444 , n9442 , n9443 );
and ( n9445 , n9444 , n6724 );
and ( n9446 , n4169 , n9115 );
or ( n9447 , n9429 , n9433 , n9437 , n9441 , n9445 , n9446 );
and ( n9448 , n9425 , n9447 );
and ( n9449 , n4169 , n3260 );
or ( n9450 , n9448 , n9449 );
and ( n9451 , n9450 , n2422 );
and ( n9452 , n4169 , n2428 );
or ( n9453 , n9451 , n9452 );
buf ( n9454 , n9453 );
buf ( n9455 , n2424 );
buf ( n9456 , n2281 );
buf ( n9457 , n2280 );
not ( n9458 , n3260 );
and ( n9459 , n7783 , n5219 );
and ( n9460 , n4159 , n9095 );
or ( n9461 , n9459 , n9460 );
and ( n9462 , n9461 , n5285 );
and ( n9463 , n7794 , n5219 );
and ( n9464 , n4159 , n9095 );
or ( n9465 , n9463 , n9464 );
and ( n9466 , n9465 , n6218 );
and ( n9467 , n7805 , n5219 );
and ( n9468 , n4159 , n9095 );
or ( n9469 , n9467 , n9468 );
and ( n9470 , n9469 , n6710 );
and ( n9471 , n5657 , n5219 );
and ( n9472 , n4159 , n9095 );
or ( n9473 , n9471 , n9472 );
and ( n9474 , n9473 , n6717 );
and ( n9475 , n7817 , n5219 );
and ( n9476 , n4159 , n9095 );
or ( n9477 , n9475 , n9476 );
and ( n9478 , n9477 , n6724 );
and ( n9479 , n4159 , n9115 );
or ( n9480 , n9462 , n9466 , n9470 , n9474 , n9478 , n9479 );
and ( n9481 , n9458 , n9480 );
and ( n9482 , n4159 , n3260 );
or ( n9483 , n9481 , n9482 );
and ( n9484 , n9483 , n2422 );
and ( n9485 , n4159 , n2428 );
or ( n9486 , n9484 , n9485 );
buf ( n9487 , n9486 );
buf ( n9488 , n2424 );
buf ( n9489 , n2281 );
buf ( n9490 , n2280 );
not ( n9491 , n3260 );
and ( n9492 , n7857 , n5219 );
and ( n9493 , n4149 , n9095 );
or ( n9494 , n9492 , n9493 );
and ( n9495 , n9494 , n5285 );
and ( n9496 , n7868 , n5219 );
and ( n9497 , n4149 , n9095 );
or ( n9498 , n9496 , n9497 );
and ( n9499 , n9498 , n6218 );
and ( n9500 , n7879 , n5219 );
and ( n9501 , n4149 , n9095 );
or ( n9502 , n9500 , n9501 );
and ( n9503 , n9502 , n6710 );
and ( n9504 , n5647 , n5219 );
and ( n9505 , n4149 , n9095 );
or ( n9506 , n9504 , n9505 );
and ( n9507 , n9506 , n6717 );
and ( n9508 , n7891 , n5219 );
and ( n9509 , n4149 , n9095 );
or ( n9510 , n9508 , n9509 );
and ( n9511 , n9510 , n6724 );
and ( n9512 , n4149 , n9115 );
or ( n9513 , n9495 , n9499 , n9503 , n9507 , n9511 , n9512 );
and ( n9514 , n9491 , n9513 );
and ( n9515 , n4149 , n3260 );
or ( n9516 , n9514 , n9515 );
and ( n9517 , n9516 , n2422 );
and ( n9518 , n4149 , n2428 );
or ( n9519 , n9517 , n9518 );
buf ( n9520 , n9519 );
buf ( n9521 , n2424 );
buf ( n9522 , n2281 );
buf ( n9523 , n2280 );
not ( n9524 , n3260 );
and ( n9525 , n7931 , n5219 );
and ( n9526 , n4139 , n9095 );
or ( n9527 , n9525 , n9526 );
and ( n9528 , n9527 , n5285 );
and ( n9529 , n7942 , n5219 );
and ( n9530 , n4139 , n9095 );
or ( n9531 , n9529 , n9530 );
and ( n9532 , n9531 , n6218 );
and ( n9533 , n7953 , n5219 );
and ( n9534 , n4139 , n9095 );
or ( n9535 , n9533 , n9534 );
and ( n9536 , n9535 , n6710 );
and ( n9537 , n5637 , n5219 );
and ( n9538 , n4139 , n9095 );
or ( n9539 , n9537 , n9538 );
and ( n9540 , n9539 , n6717 );
and ( n9541 , n7965 , n5219 );
and ( n9542 , n4139 , n9095 );
or ( n9543 , n9541 , n9542 );
and ( n9544 , n9543 , n6724 );
and ( n9545 , n4139 , n9115 );
or ( n9546 , n9528 , n9532 , n9536 , n9540 , n9544 , n9545 );
and ( n9547 , n9524 , n9546 );
and ( n9548 , n4139 , n3260 );
or ( n9549 , n9547 , n9548 );
and ( n9550 , n9549 , n2422 );
and ( n9551 , n4139 , n2428 );
or ( n9552 , n9550 , n9551 );
buf ( n9553 , n9552 );
buf ( n9554 , n2424 );
buf ( n9555 , n2281 );
buf ( n9556 , n2280 );
not ( n9557 , n3260 );
and ( n9558 , n8005 , n5219 );
and ( n9559 , n4129 , n9095 );
or ( n9560 , n9558 , n9559 );
and ( n9561 , n9560 , n5285 );
and ( n9562 , n8016 , n5219 );
and ( n9563 , n4129 , n9095 );
or ( n9564 , n9562 , n9563 );
and ( n9565 , n9564 , n6218 );
and ( n9566 , n8027 , n5219 );
and ( n9567 , n4129 , n9095 );
or ( n9568 , n9566 , n9567 );
and ( n9569 , n9568 , n6710 );
and ( n9570 , n5627 , n5219 );
and ( n9571 , n4129 , n9095 );
or ( n9572 , n9570 , n9571 );
and ( n9573 , n9572 , n6717 );
and ( n9574 , n8039 , n5219 );
and ( n9575 , n4129 , n9095 );
or ( n9576 , n9574 , n9575 );
and ( n9577 , n9576 , n6724 );
and ( n9578 , n4129 , n9115 );
or ( n9579 , n9561 , n9565 , n9569 , n9573 , n9577 , n9578 );
and ( n9580 , n9557 , n9579 );
and ( n9581 , n4129 , n3260 );
or ( n9582 , n9580 , n9581 );
and ( n9583 , n9582 , n2422 );
and ( n9584 , n4129 , n2428 );
xor ( n9585 , n9583 , n9584 );
buf ( n9586 , n9585 );
buf ( n9587 , n2424 );
buf ( n9588 , n2281 );
buf ( n9589 , n2280 );
not ( n9590 , n3260 );
and ( n9591 , n8079 , n5219 );
and ( n9592 , n4119 , n9095 );
or ( n9593 , n9591 , n9592 );
and ( n9594 , n9593 , n5285 );
and ( n9595 , n8090 , n5219 );
and ( n9596 , n4119 , n9095 );
or ( n9597 , n9595 , n9596 );
and ( n9598 , n9597 , n6218 );
and ( n9599 , n8101 , n5219 );
and ( n9600 , n4119 , n9095 );
or ( n9601 , n9599 , n9600 );
and ( n9602 , n9601 , n6710 );
and ( n9603 , n5617 , n5219 );
and ( n9604 , n4119 , n9095 );
or ( n9605 , n9603 , n9604 );
and ( n9606 , n9605 , n6717 );
and ( n9607 , n8113 , n5219 );
and ( n9608 , n4119 , n9095 );
or ( n9609 , n9607 , n9608 );
and ( n9610 , n9609 , n6724 );
and ( n9611 , n4119 , n9115 );
or ( n9612 , n9594 , n9598 , n9602 , n9606 , n9610 , n9611 );
and ( n9613 , n9590 , n9612 );
and ( n9614 , n4119 , n3260 );
or ( n9615 , n9613 , n9614 );
and ( n9616 , n9615 , n2422 );
and ( n9617 , n4119 , n2428 );
or ( n9618 , n9616 , n9617 );
buf ( n9619 , n9618 );
buf ( n9620 , n2424 );
buf ( n9621 , n2281 );
buf ( n9622 , n2280 );
not ( n9623 , n3260 );
and ( n9624 , n8153 , n5219 );
and ( n9625 , n4109 , n9095 );
or ( n9626 , n9624 , n9625 );
and ( n9627 , n9626 , n5285 );
and ( n9628 , n8164 , n5219 );
and ( n9629 , n4109 , n9095 );
or ( n9630 , n9628 , n9629 );
and ( n9631 , n9630 , n6218 );
and ( n9632 , n8175 , n5219 );
and ( n9633 , n4109 , n9095 );
or ( n9634 , n9632 , n9633 );
and ( n9635 , n9634 , n6710 );
and ( n9636 , n5607 , n5219 );
and ( n9637 , n4109 , n9095 );
or ( n9638 , n9636 , n9637 );
and ( n9639 , n9638 , n6717 );
and ( n9640 , n8187 , n5219 );
and ( n9641 , n4109 , n9095 );
or ( n9642 , n9640 , n9641 );
and ( n9643 , n9642 , n6724 );
and ( n9644 , n4109 , n9115 );
or ( n9645 , n9627 , n9631 , n9635 , n9639 , n9643 , n9644 );
and ( n9646 , n9623 , n9645 );
and ( n9647 , n4109 , n3260 );
or ( n9648 , n9646 , n9647 );
and ( n9649 , n9648 , n2422 );
and ( n9650 , n4109 , n2428 );
or ( n9651 , n9649 , n9650 );
buf ( n9652 , n9651 );
buf ( n9653 , n2424 );
buf ( n9654 , n2281 );
buf ( n9655 , n2280 );
not ( n9656 , n3260 );
and ( n9657 , n8227 , n5219 );
and ( n9658 , n4099 , n9095 );
or ( n9659 , n9657 , n9658 );
and ( n9660 , n9659 , n5285 );
and ( n9661 , n8238 , n5219 );
and ( n9662 , n4099 , n9095 );
or ( n9663 , n9661 , n9662 );
and ( n9664 , n9663 , n6218 );
and ( n9665 , n8249 , n5219 );
and ( n9666 , n4099 , n9095 );
or ( n9667 , n9665 , n9666 );
and ( n9668 , n9667 , n6710 );
and ( n9669 , n5597 , n5219 );
and ( n9670 , n4099 , n9095 );
or ( n9671 , n9669 , n9670 );
and ( n9672 , n9671 , n6717 );
and ( n9673 , n8261 , n5219 );
and ( n9674 , n4099 , n9095 );
or ( n9675 , n9673 , n9674 );
and ( n9676 , n9675 , n6724 );
and ( n9677 , n4099 , n9115 );
or ( n9678 , n9660 , n9664 , n9668 , n9672 , n9676 , n9677 );
and ( n9679 , n9656 , n9678 );
and ( n9680 , n4099 , n3260 );
or ( n9681 , n9679 , n9680 );
and ( n9682 , n9681 , n2422 );
and ( n9683 , n4099 , n2428 );
or ( n9684 , n9682 , n9683 );
buf ( n9685 , n9684 );
buf ( n9686 , n2424 );
buf ( n9687 , n2281 );
buf ( n9688 , n2280 );
not ( n9689 , n3260 );
and ( n9690 , n8301 , n5219 );
and ( n9691 , n4089 , n9095 );
or ( n9692 , n9690 , n9691 );
and ( n9693 , n9692 , n5285 );
and ( n9694 , n8312 , n5219 );
and ( n9695 , n4089 , n9095 );
or ( n9696 , n9694 , n9695 );
and ( n9697 , n9696 , n6218 );
and ( n9698 , n8323 , n5219 );
and ( n9699 , n4089 , n9095 );
or ( n9700 , n9698 , n9699 );
and ( n9701 , n9700 , n6710 );
and ( n9702 , n5587 , n5219 );
and ( n9703 , n4089 , n9095 );
or ( n9704 , n9702 , n9703 );
and ( n9705 , n9704 , n6717 );
and ( n9706 , n8335 , n5219 );
and ( n9707 , n4089 , n9095 );
or ( n9708 , n9706 , n9707 );
and ( n9709 , n9708 , n6724 );
and ( n9710 , n4089 , n9115 );
or ( n9711 , n9693 , n9697 , n9701 , n9705 , n9709 , n9710 );
and ( n9712 , n9689 , n9711 );
and ( n9713 , n4089 , n3260 );
or ( n9714 , n9712 , n9713 );
and ( n9715 , n9714 , n2422 );
and ( n9716 , n4089 , n2428 );
or ( n9717 , n9715 , n9716 );
buf ( n9718 , n9717 );
buf ( n9719 , n2424 );
buf ( n9720 , n2281 );
buf ( n9721 , n2280 );
not ( n9722 , n3260 );
and ( n9723 , n8375 , n5219 );
and ( n9724 , n4079 , n9095 );
or ( n9725 , n9723 , n9724 );
and ( n9726 , n9725 , n5285 );
and ( n9727 , n8386 , n5219 );
and ( n9728 , n4079 , n9095 );
or ( n9729 , n9727 , n9728 );
and ( n9730 , n9729 , n6218 );
and ( n9731 , n8397 , n5219 );
and ( n9732 , n4079 , n9095 );
or ( n9733 , n9731 , n9732 );
and ( n9734 , n9733 , n6710 );
and ( n9735 , n5577 , n5219 );
and ( n9736 , n4079 , n9095 );
or ( n9737 , n9735 , n9736 );
and ( n9738 , n9737 , n6717 );
and ( n9739 , n8409 , n5219 );
and ( n9740 , n4079 , n9095 );
or ( n9741 , n9739 , n9740 );
and ( n9742 , n9741 , n6724 );
and ( n9743 , n4079 , n9115 );
or ( n9744 , n9726 , n9730 , n9734 , n9738 , n9742 , n9743 );
and ( n9745 , n9722 , n9744 );
and ( n9746 , n4079 , n3260 );
or ( n9747 , n9745 , n9746 );
and ( n9748 , n9747 , n2422 );
and ( n9749 , n4079 , n2428 );
or ( n9750 , n9748 , n9749 );
buf ( n9751 , n9750 );
buf ( n9752 , n2424 );
buf ( n9753 , n2281 );
buf ( n9754 , n2280 );
not ( n9755 , n3260 );
and ( n9756 , n8449 , n5219 );
and ( n9757 , n4069 , n9095 );
or ( n9758 , n9756 , n9757 );
and ( n9759 , n9758 , n5285 );
and ( n9760 , n8460 , n5219 );
and ( n9761 , n4069 , n9095 );
or ( n9762 , n9760 , n9761 );
and ( n9763 , n9762 , n6218 );
and ( n9764 , n8471 , n5219 );
and ( n9765 , n4069 , n9095 );
or ( n9766 , n9764 , n9765 );
and ( n9767 , n9766 , n6710 );
and ( n9768 , n5529 , n5219 );
and ( n9769 , n4069 , n9095 );
or ( n9770 , n9768 , n9769 );
and ( n9771 , n9770 , n6717 );
and ( n9772 , n8483 , n5219 );
and ( n9773 , n4069 , n9095 );
or ( n9774 , n9772 , n9773 );
and ( n9775 , n9774 , n6724 );
and ( n9776 , n4069 , n9115 );
or ( n9777 , n9759 , n9763 , n9767 , n9771 , n9775 , n9776 );
and ( n9778 , n9755 , n9777 );
and ( n9779 , n4069 , n3260 );
or ( n9780 , n9778 , n9779 );
and ( n9781 , n9780 , n2422 );
and ( n9782 , n4069 , n2428 );
or ( n9783 , n9781 , n9782 );
buf ( n9784 , n9783 );
buf ( n9785 , n2424 );
buf ( n9786 , n2281 );
buf ( n9787 , n2280 );
not ( n9788 , n3260 );
and ( n9789 , n8523 , n5219 );
and ( n9790 , n4059 , n9095 );
or ( n9791 , n9789 , n9790 );
and ( n9792 , n9791 , n5285 );
and ( n9793 , n8534 , n5219 );
and ( n9794 , n4059 , n9095 );
or ( n9795 , n9793 , n9794 );
and ( n9796 , n9795 , n6218 );
and ( n9797 , n8545 , n5219 );
and ( n9798 , n4059 , n9095 );
or ( n9799 , n9797 , n9798 );
and ( n9800 , n9799 , n6710 );
and ( n9801 , n5526 , n5219 );
and ( n9802 , n4059 , n9095 );
or ( n9803 , n9801 , n9802 );
and ( n9804 , n9803 , n6717 );
and ( n9805 , n8557 , n5219 );
and ( n9806 , n4059 , n9095 );
or ( n9807 , n9805 , n9806 );
and ( n9808 , n9807 , n6724 );
and ( n9809 , n4059 , n9115 );
or ( n9810 , n9792 , n9796 , n9800 , n9804 , n9808 , n9809 );
and ( n9811 , n9788 , n9810 );
and ( n9812 , n4059 , n3260 );
or ( n9813 , n9811 , n9812 );
and ( n9814 , n9813 , n2422 );
and ( n9815 , n4059 , n2428 );
or ( n9816 , n9814 , n9815 );
buf ( n9817 , n9816 );
buf ( n9818 , n2424 );
buf ( n9819 , n2281 );
buf ( n9820 , n2280 );
not ( n9821 , n3260 );
and ( n9822 , n8597 , n5219 );
and ( n9823 , n4049 , n9095 );
or ( n9824 , n9822 , n9823 );
and ( n9825 , n9824 , n5285 );
and ( n9826 , n8608 , n5219 );
and ( n9827 , n4049 , n9095 );
or ( n9828 , n9826 , n9827 );
and ( n9829 , n9828 , n6218 );
and ( n9830 , n8619 , n5219 );
and ( n9831 , n4049 , n9095 );
or ( n9832 , n9830 , n9831 );
and ( n9833 , n9832 , n6710 );
and ( n9834 , n5523 , n5219 );
and ( n9835 , n4049 , n9095 );
or ( n9836 , n9834 , n9835 );
and ( n9837 , n9836 , n6717 );
and ( n9838 , n8631 , n5219 );
and ( n9839 , n4049 , n9095 );
or ( n9840 , n9838 , n9839 );
and ( n9841 , n9840 , n6724 );
and ( n9842 , n4049 , n9115 );
or ( n9843 , n9825 , n9829 , n9833 , n9837 , n9841 , n9842 );
and ( n9844 , n9821 , n9843 );
and ( n9845 , n4049 , n3260 );
or ( n9846 , n9844 , n9845 );
and ( n9847 , n9846 , n2422 );
and ( n9848 , n4049 , n2428 );
or ( n9849 , n9847 , n9848 );
buf ( n9850 , n9849 );
buf ( n9851 , n2424 );
buf ( n9852 , n2281 );
buf ( n9853 , n2280 );
not ( n9854 , n3260 );
and ( n9855 , n8671 , n5219 );
and ( n9856 , n4039 , n9095 );
or ( n9857 , n9855 , n9856 );
and ( n9858 , n9857 , n5285 );
and ( n9859 , n8682 , n5219 );
and ( n9860 , n4039 , n9095 );
or ( n9861 , n9859 , n9860 );
and ( n9862 , n9861 , n6218 );
and ( n9863 , n8693 , n5219 );
and ( n9864 , n4039 , n9095 );
or ( n9865 , n9863 , n9864 );
and ( n9866 , n9865 , n6710 );
and ( n9867 , n5520 , n5219 );
and ( n9868 , n4039 , n9095 );
or ( n9869 , n9867 , n9868 );
and ( n9870 , n9869 , n6717 );
and ( n9871 , n8705 , n5219 );
and ( n9872 , n4039 , n9095 );
or ( n9873 , n9871 , n9872 );
and ( n9874 , n9873 , n6724 );
and ( n9875 , n4039 , n9115 );
or ( n9876 , n9858 , n9862 , n9866 , n9870 , n9874 , n9875 );
and ( n9877 , n9854 , n9876 );
and ( n9878 , n4039 , n3260 );
or ( n9879 , n9877 , n9878 );
and ( n9880 , n9879 , n2422 );
and ( n9881 , n4039 , n2428 );
or ( n9882 , n9880 , n9881 );
buf ( n9883 , n9882 );
buf ( n9884 , n2424 );
buf ( n9885 , n2281 );
buf ( n9886 , n2280 );
not ( n9887 , n3260 );
and ( n9888 , n8745 , n5219 );
and ( n9889 , n4029 , n9095 );
or ( n9890 , n9888 , n9889 );
and ( n9891 , n9890 , n5285 );
and ( n9892 , n8756 , n5219 );
and ( n9893 , n4029 , n9095 );
or ( n9894 , n9892 , n9893 );
and ( n9895 , n9894 , n6218 );
and ( n9896 , n8767 , n5219 );
and ( n9897 , n4029 , n9095 );
or ( n9898 , n9896 , n9897 );
and ( n9899 , n9898 , n6710 );
and ( n9900 , n5517 , n5219 );
and ( n9901 , n4029 , n9095 );
or ( n9902 , n9900 , n9901 );
and ( n9903 , n9902 , n6717 );
and ( n9904 , n8779 , n5219 );
and ( n9905 , n4029 , n9095 );
or ( n9906 , n9904 , n9905 );
and ( n9907 , n9906 , n6724 );
and ( n9908 , n4029 , n9115 );
or ( n9909 , n9891 , n9895 , n9899 , n9903 , n9907 , n9908 );
and ( n9910 , n9887 , n9909 );
and ( n9911 , n4029 , n3260 );
or ( n9912 , n9910 , n9911 );
and ( n9913 , n9912 , n2422 );
and ( n9914 , n4029 , n2428 );
or ( n9915 , n9913 , n9914 );
buf ( n9916 , n9915 );
buf ( n9917 , n2424 );
buf ( n9918 , n2281 );
buf ( n9919 , n2280 );
not ( n9920 , n3260 );
and ( n9921 , n8819 , n5219 );
and ( n9922 , n4019 , n9095 );
or ( n9923 , n9921 , n9922 );
and ( n9924 , n9923 , n5285 );
and ( n9925 , n8830 , n5219 );
and ( n9926 , n4019 , n9095 );
or ( n9927 , n9925 , n9926 );
and ( n9928 , n9927 , n6218 );
and ( n9929 , n8841 , n5219 );
and ( n9930 , n4019 , n9095 );
or ( n9931 , n9929 , n9930 );
and ( n9932 , n9931 , n6710 );
and ( n9933 , n5514 , n5219 );
and ( n9934 , n4019 , n9095 );
or ( n9935 , n9933 , n9934 );
and ( n9936 , n9935 , n6717 );
and ( n9937 , n8853 , n5219 );
and ( n9938 , n4019 , n9095 );
or ( n9939 , n9937 , n9938 );
and ( n9940 , n9939 , n6724 );
and ( n9941 , n4019 , n9115 );
or ( n9942 , n9924 , n9928 , n9932 , n9936 , n9940 , n9941 );
and ( n9943 , n9920 , n9942 );
and ( n9944 , n4019 , n3260 );
or ( n9945 , n9943 , n9944 );
and ( n9946 , n9945 , n2422 );
and ( n9947 , n4019 , n2428 );
or ( n9948 , n9946 , n9947 );
buf ( n9949 , n9948 );
buf ( n9950 , n2424 );
buf ( n9951 , n2281 );
buf ( n9952 , n2280 );
not ( n9953 , n3260 );
and ( n9954 , n8893 , n5219 );
and ( n9955 , n4009 , n9095 );
or ( n9956 , n9954 , n9955 );
and ( n9957 , n9956 , n5285 );
and ( n9958 , n8904 , n5219 );
and ( n9959 , n4009 , n9095 );
or ( n9960 , n9958 , n9959 );
and ( n9961 , n9960 , n6218 );
and ( n9962 , n8915 , n5219 );
and ( n9963 , n4009 , n9095 );
or ( n9964 , n9962 , n9963 );
and ( n9965 , n9964 , n6710 );
and ( n9966 , n5511 , n5219 );
and ( n9967 , n4009 , n9095 );
or ( n9968 , n9966 , n9967 );
and ( n9969 , n9968 , n6717 );
and ( n9970 , n8927 , n5219 );
and ( n9971 , n4009 , n9095 );
or ( n9972 , n9970 , n9971 );
and ( n9973 , n9972 , n6724 );
and ( n9974 , n4009 , n9115 );
or ( n9975 , n9957 , n9961 , n9965 , n9969 , n9973 , n9974 );
and ( n9976 , n9953 , n9975 );
and ( n9977 , n4009 , n3260 );
or ( n9978 , n9976 , n9977 );
and ( n9979 , n9978 , n2422 );
and ( n9980 , n4009 , n2428 );
or ( n9981 , n9979 , n9980 );
buf ( n9982 , n9981 );
buf ( n9983 , n2424 );
buf ( n9984 , n2281 );
buf ( n9985 , n2280 );
not ( n9986 , n3260 );
and ( n9987 , n8967 , n5219 );
and ( n9988 , n3999 , n9095 );
or ( n9989 , n9987 , n9988 );
and ( n9990 , n9989 , n5285 );
and ( n9991 , n8978 , n5219 );
and ( n9992 , n3999 , n9095 );
or ( n9993 , n9991 , n9992 );
and ( n9994 , n9993 , n6218 );
and ( n9995 , n8989 , n5219 );
and ( n9996 , n3999 , n9095 );
or ( n9997 , n9995 , n9996 );
and ( n9998 , n9997 , n6710 );
and ( n9999 , n5508 , n5219 );
and ( n10000 , n3999 , n9095 );
or ( n10001 , n9999 , n10000 );
and ( n10002 , n10001 , n6717 );
and ( n10003 , n9001 , n5219 );
and ( n10004 , n3999 , n9095 );
or ( n10005 , n10003 , n10004 );
and ( n10006 , n10005 , n6724 );
and ( n10007 , n3999 , n9115 );
or ( n10008 , n9990 , n9994 , n9998 , n10002 , n10006 , n10007 );
and ( n10009 , n9986 , n10008 );
and ( n10010 , n3999 , n3260 );
or ( n10011 , n10009 , n10010 );
and ( n10012 , n10011 , n2422 );
and ( n10013 , n3999 , n2428 );
or ( n10014 , n10012 , n10013 );
buf ( n10015 , n10014 );
buf ( n10016 , n2424 );
buf ( n10017 , n2281 );
buf ( n10018 , n2280 );
not ( n10019 , n3260 );
and ( n10020 , n9041 , n5219 );
and ( n10021 , n3989 , n9095 );
or ( n10022 , n10020 , n10021 );
and ( n10023 , n10022 , n5285 );
and ( n10024 , n9052 , n5219 );
and ( n10025 , n3989 , n9095 );
or ( n10026 , n10024 , n10025 );
and ( n10027 , n10026 , n6218 );
and ( n10028 , n9063 , n5219 );
and ( n10029 , n3989 , n9095 );
or ( n10030 , n10028 , n10029 );
and ( n10031 , n10030 , n6710 );
and ( n10032 , n5505 , n5219 );
and ( n10033 , n3989 , n9095 );
or ( n10034 , n10032 , n10033 );
and ( n10035 , n10034 , n6717 );
and ( n10036 , n9075 , n5219 );
and ( n10037 , n3989 , n9095 );
or ( n10038 , n10036 , n10037 );
and ( n10039 , n10038 , n6724 );
and ( n10040 , n3989 , n9115 );
or ( n10041 , n10023 , n10027 , n10031 , n10035 , n10039 , n10040 );
and ( n10042 , n10019 , n10041 );
and ( n10043 , n3989 , n3260 );
or ( n10044 , n10042 , n10043 );
and ( n10045 , n10044 , n2422 );
and ( n10046 , n3989 , n2428 );
or ( n10047 , n10045 , n10046 );
buf ( n10048 , n10047 );
buf ( n10049 , n2424 );
buf ( n10050 , n2281 );
buf ( n10051 , n2280 );
not ( n10052 , n3260 );
not ( n10053 , n7021 );
and ( n10054 , n10053 , n7019 );
xor ( n10055 , n7019 , n3770 );
and ( n10056 , n9021 , n9022 );
xor ( n10057 , n10055 , n10056 );
and ( n10058 , n10057 , n7021 );
or ( n10059 , n10054 , n10058 );
and ( n10060 , n10059 , n5289 );
and ( n10061 , n10059 , n5287 );
not ( n10062 , n3290 );
not ( n10063 , n3770 );
and ( n10064 , n10063 , n4301 );
xor ( n10065 , n4302 , n4573 );
and ( n10066 , n10065 , n3770 );
or ( n10067 , n10064 , n10066 );
and ( n10068 , n10062 , n10067 );
not ( n10069 , n4999 );
and ( n10070 , n10069 , n2424 );
and ( n10071 , n9032 , n9033 );
and ( n10072 , n10071 , n4999 );
or ( n10073 , n10070 , n10072 );
and ( n10074 , n10073 , n3290 );
or ( n10075 , n10068 , n10074 );
and ( n10076 , n10075 , n5152 );
and ( n10077 , n10067 , n5154 );
or ( n10078 , n10060 , n10061 , n10076 , n10077 );
and ( n10079 , n10078 , n5219 );
and ( n10080 , n3979 , n9095 );
or ( n10081 , n10079 , n10080 );
and ( n10082 , n10081 , n5285 );
not ( n10083 , n6201 );
and ( n10084 , n10083 , n6199 );
xor ( n10085 , n6199 , n5852 );
and ( n10086 , n9048 , n9049 );
xor ( n10087 , n10085 , n10086 );
and ( n10088 , n10087 , n6201 );
or ( n10089 , n10084 , n10088 );
and ( n10090 , n10089 , n5219 );
and ( n10091 , n3979 , n9095 );
or ( n10092 , n10090 , n10091 );
and ( n10093 , n10092 , n6218 );
not ( n10094 , n6694 );
and ( n10095 , n10094 , n6692 );
xor ( n10096 , n6692 , n6345 );
and ( n10097 , n9059 , n9060 );
xor ( n10098 , n10096 , n10097 );
and ( n10099 , n10098 , n6694 );
or ( n10100 , n10095 , n10099 );
and ( n10101 , n10100 , n5219 );
and ( n10102 , n3979 , n9095 );
or ( n10103 , n10101 , n10102 );
and ( n10104 , n10103 , n6710 );
and ( n10105 , n5502 , n5219 );
and ( n10106 , n3979 , n9095 );
or ( n10107 , n10105 , n10106 );
and ( n10108 , n10107 , n6717 );
not ( n10109 , n5502 );
and ( n10110 , n9073 , n9074 );
xor ( n10111 , n10109 , n10110 );
and ( n10112 , n10111 , n5219 );
and ( n10113 , n3979 , n9095 );
or ( n10114 , n10112 , n10113 );
and ( n10115 , n10114 , n6724 );
and ( n10116 , n3979 , n9115 );
or ( n10117 , n10082 , n10093 , n10104 , n10108 , n10115 , n10116 );
and ( n10118 , n10052 , n10117 );
and ( n10119 , n3979 , n3260 );
or ( n10120 , n10118 , n10119 );
and ( n10121 , n10120 , n2422 );
and ( n10122 , n3979 , n2428 );
or ( n10123 , n10121 , n10122 );
buf ( n10124 , n10123 );
buf ( n10125 , n2424 );
buf ( n10126 , n2281 );
buf ( n10127 , n2280 );
not ( n10128 , n3260 );
not ( n10129 , n7021 );
and ( n10130 , n10129 , n2424 );
and ( n10131 , n10055 , n10056 );
and ( n10132 , n10131 , n7021 );
or ( n10133 , n10130 , n10132 );
and ( n10134 , n10133 , n5289 );
and ( n10135 , n10133 , n5287 );
not ( n10136 , n3290 );
not ( n10137 , n3770 );
and ( n10138 , n10137 , n4293 );
xor ( n10139 , n4294 , n4574 );
and ( n10140 , n10139 , n3770 );
or ( n10141 , n10138 , n10140 );
and ( n10142 , n10136 , n10141 );
and ( n10143 , n2424 , n3290 );
or ( n10144 , n10142 , n10143 );
and ( n10145 , n10144 , n5152 );
and ( n10146 , n10141 , n5154 );
or ( n10147 , n10134 , n10135 , n10145 , n10146 );
and ( n10148 , n10147 , n5219 );
and ( n10149 , n3815 , n9095 );
or ( n10150 , n10148 , n10149 );
and ( n10151 , n10150 , n5285 );
not ( n10152 , n6201 );
and ( n10153 , n10152 , n2424 );
and ( n10154 , n10085 , n10086 );
and ( n10155 , n10154 , n6201 );
or ( n10156 , n10153 , n10155 );
and ( n10157 , n10156 , n5219 );
and ( n10158 , n3815 , n9095 );
or ( n10159 , n10157 , n10158 );
and ( n10160 , n10159 , n6218 );
not ( n10161 , n6694 );
and ( n10162 , n10161 , n2424 );
and ( n10163 , n10096 , n10097 );
and ( n10164 , n10163 , n6694 );
or ( n10165 , n10162 , n10164 );
and ( n10166 , n10165 , n5219 );
and ( n10167 , n3815 , n9095 );
or ( n10168 , n10166 , n10167 );
and ( n10169 , n10168 , n6710 );
and ( n10170 , n5499 , n5219 );
and ( n10171 , n3815 , n9095 );
or ( n10172 , n10170 , n10171 );
and ( n10173 , n10172 , n6717 );
not ( n10174 , n5499 );
and ( n10175 , n10109 , n10110 );
xor ( n10176 , n10174 , n10175 );
and ( n10177 , n10176 , n5219 );
and ( n10178 , n3815 , n9095 );
or ( n10179 , n10177 , n10178 );
and ( n10180 , n10179 , n6724 );
and ( n10181 , n3815 , n9115 );
or ( n10182 , n10151 , n10160 , n10169 , n10173 , n10180 , n10181 );
and ( n10183 , n10128 , n10182 );
and ( n10184 , n3815 , n3260 );
or ( n10185 , n10183 , n10184 );
and ( n10186 , n10185 , n2422 );
and ( n10187 , n3815 , n2428 );
or ( n10188 , n10186 , n10187 );
buf ( n10189 , n10188 );
buf ( n10190 , n2424 );
buf ( n10191 , n2281 );
buf ( n10192 , n2280 );
not ( n10193 , n3260 );
buf ( n10194 , n2424 );
not ( n10195 , n3290 );
and ( n10196 , n10195 , n4578 );
and ( n10197 , n2424 , n3290 );
or ( n10198 , n10196 , n10197 );
and ( n10199 , n10198 , n5152 );
and ( n10200 , n4578 , n5154 );
or ( n10201 , n2424 , n10194 , n10199 , n10200 );
and ( n10202 , n10201 , n5219 );
and ( n10203 , n3764 , n9095 );
or ( n10204 , n10202 , n10203 );
and ( n10205 , n10204 , n5285 );
and ( n10206 , n3764 , n9095 );
and ( n10207 , n10206 , n6218 );
and ( n10208 , n3764 , n9095 );
and ( n10209 , n10208 , n6710 );
and ( n10210 , n5496 , n5219 );
and ( n10211 , n3764 , n9095 );
or ( n10212 , n10210 , n10211 );
and ( n10213 , n10212 , n6717 );
not ( n10214 , n5496 );
and ( n10215 , n10174 , n10175 );
xor ( n10216 , n10214 , n10215 );
and ( n10217 , n10216 , n5219 );
and ( n10218 , n3764 , n9095 );
or ( n10219 , n10217 , n10218 );
and ( n10220 , n10219 , n6724 );
and ( n10221 , n3764 , n9115 );
or ( n10222 , n10205 , n10207 , n10209 , n10213 , n10220 , n10221 );
and ( n10223 , n10193 , n10222 );
and ( n10224 , n3764 , n3260 );
or ( n10225 , n10223 , n10224 );
and ( n10226 , n10225 , n2422 );
and ( n10227 , n3764 , n2428 );
or ( n10228 , n10226 , n10227 );
buf ( n10229 , n10228 );
buf ( n10230 , n2424 );
buf ( n10231 , n2281 );
buf ( n10232 , n2280 );
not ( n10233 , n3260 );
and ( n10234 , n5156 , n5249 );
or ( n10235 , n5219 , n5280 );
or ( n10236 , n10235 , n5188 );
buf ( n10237 , n10236 );
and ( n10238 , n3793 , n10237 );
or ( n10239 , n10234 , n10238 );
and ( n10240 , n10239 , n5285 );
and ( n10241 , n6207 , n5249 );
and ( n10242 , n3793 , n10237 );
or ( n10243 , n10241 , n10242 );
and ( n10244 , n10243 , n6218 );
and ( n10245 , n6700 , n5249 );
and ( n10246 , n3793 , n10237 );
or ( n10247 , n10245 , n10246 );
and ( n10248 , n10247 , n6710 );
and ( n10249 , n5492 , n5249 );
and ( n10250 , n3793 , n10237 );
or ( n10251 , n10249 , n10250 );
and ( n10252 , n10251 , n6717 );
and ( n10253 , n5492 , n5249 );
and ( n10254 , n3793 , n10237 );
or ( n10255 , n10253 , n10254 );
and ( n10256 , n10255 , n6724 );
and ( n10257 , n3793 , n9115 );
or ( n10258 , n10240 , n10244 , n10248 , n10252 , n10256 , n10257 );
and ( n10259 , n10233 , n10258 );
and ( n10260 , n3793 , n3260 );
or ( n10261 , n10259 , n10260 );
and ( n10262 , n10261 , n2422 );
and ( n10263 , n3793 , n2428 );
or ( n10264 , n10262 , n10263 );
buf ( n10265 , n10264 );
buf ( n10266 , n2424 );
buf ( n10267 , n2281 );
buf ( n10268 , n2280 );
not ( n10269 , n3260 );
and ( n10270 , n7043 , n5249 );
and ( n10271 , n3783 , n10237 );
or ( n10272 , n10270 , n10271 );
and ( n10273 , n10272 , n5285 );
and ( n10274 , n7054 , n5249 );
and ( n10275 , n3783 , n10237 );
or ( n10276 , n10274 , n10275 );
and ( n10277 , n10276 , n6218 );
and ( n10278 , n7065 , n5249 );
and ( n10279 , n3783 , n10237 );
or ( n10280 , n10278 , n10279 );
and ( n10281 , n10280 , n6710 );
and ( n10282 , n5757 , n5249 );
and ( n10283 , n3783 , n10237 );
or ( n10284 , n10282 , n10283 );
and ( n10285 , n10284 , n6717 );
and ( n10286 , n7077 , n5249 );
and ( n10287 , n3783 , n10237 );
or ( n10288 , n10286 , n10287 );
and ( n10289 , n10288 , n6724 );
and ( n10290 , n3783 , n9115 );
or ( n10291 , n10273 , n10277 , n10281 , n10285 , n10289 , n10290 );
and ( n10292 , n10269 , n10291 );
and ( n10293 , n3783 , n3260 );
or ( n10294 , n10292 , n10293 );
and ( n10295 , n10294 , n2422 );
and ( n10296 , n3783 , n2428 );
or ( n10297 , n10295 , n10296 );
buf ( n10298 , n10297 );
buf ( n10299 , n2424 );
buf ( n10300 , n2281 );
buf ( n10301 , n2280 );
not ( n10302 , n3260 );
and ( n10303 , n7117 , n5249 );
and ( n10304 , n4255 , n10237 );
or ( n10305 , n10303 , n10304 );
and ( n10306 , n10305 , n5285 );
and ( n10307 , n7128 , n5249 );
and ( n10308 , n4255 , n10237 );
or ( n10309 , n10307 , n10308 );
and ( n10310 , n10309 , n6218 );
and ( n10311 , n7139 , n5249 );
and ( n10312 , n4255 , n10237 );
or ( n10313 , n10311 , n10312 );
and ( n10314 , n10313 , n6710 );
and ( n10315 , n5747 , n5249 );
and ( n10316 , n4255 , n10237 );
or ( n10317 , n10315 , n10316 );
and ( n10318 , n10317 , n6717 );
and ( n10319 , n7151 , n5249 );
and ( n10320 , n4255 , n10237 );
or ( n10321 , n10319 , n10320 );
and ( n10322 , n10321 , n6724 );
and ( n10323 , n4255 , n9115 );
or ( n10324 , n10306 , n10310 , n10314 , n10318 , n10322 , n10323 );
and ( n10325 , n10302 , n10324 );
and ( n10326 , n4255 , n3260 );
or ( n10327 , n10325 , n10326 );
and ( n10328 , n10327 , n2422 );
and ( n10329 , n4255 , n2428 );
or ( n10330 , n10328 , n10329 );
buf ( n10331 , n10330 );
buf ( n10332 , n2424 );
buf ( n10333 , n2281 );
buf ( n10334 , n2280 );
not ( n10335 , n3260 );
and ( n10336 , n7191 , n5249 );
and ( n10337 , n4241 , n10237 );
or ( n10338 , n10336 , n10337 );
and ( n10339 , n10338 , n5285 );
and ( n10340 , n7202 , n5249 );
and ( n10341 , n4241 , n10237 );
or ( n10342 , n10340 , n10341 );
and ( n10343 , n10342 , n6218 );
and ( n10344 , n7213 , n5249 );
and ( n10345 , n4241 , n10237 );
or ( n10346 , n10344 , n10345 );
and ( n10347 , n10346 , n6710 );
and ( n10348 , n5737 , n5249 );
and ( n10349 , n4241 , n10237 );
or ( n10350 , n10348 , n10349 );
and ( n10351 , n10350 , n6717 );
and ( n10352 , n7225 , n5249 );
and ( n10353 , n4241 , n10237 );
or ( n10354 , n10352 , n10353 );
and ( n10355 , n10354 , n6724 );
and ( n10356 , n4241 , n9115 );
or ( n10357 , n10339 , n10343 , n10347 , n10351 , n10355 , n10356 );
and ( n10358 , n10335 , n10357 );
and ( n10359 , n4241 , n3260 );
or ( n10360 , n10358 , n10359 );
and ( n10361 , n10360 , n2422 );
and ( n10362 , n4241 , n2428 );
or ( n10363 , n10361 , n10362 );
buf ( n10364 , n10363 );
buf ( n10365 , n2424 );
buf ( n10366 , n2281 );
buf ( n10367 , n2280 );
not ( n10368 , n3260 );
and ( n10369 , n7265 , n5249 );
and ( n10370 , n4231 , n10237 );
or ( n10371 , n10369 , n10370 );
and ( n10372 , n10371 , n5285 );
and ( n10373 , n7276 , n5249 );
and ( n10374 , n4231 , n10237 );
or ( n10375 , n10373 , n10374 );
and ( n10376 , n10375 , n6218 );
and ( n10377 , n7287 , n5249 );
and ( n10378 , n4231 , n10237 );
or ( n10379 , n10377 , n10378 );
and ( n10380 , n10379 , n6710 );
and ( n10381 , n5727 , n5249 );
and ( n10382 , n4231 , n10237 );
or ( n10383 , n10381 , n10382 );
and ( n10384 , n10383 , n6717 );
and ( n10385 , n7299 , n5249 );
and ( n10386 , n4231 , n10237 );
or ( n10387 , n10385 , n10386 );
and ( n10388 , n10387 , n6724 );
and ( n10389 , n4231 , n9115 );
or ( n10390 , n10372 , n10376 , n10380 , n10384 , n10388 , n10389 );
and ( n10391 , n10368 , n10390 );
and ( n10392 , n4231 , n3260 );
or ( n10393 , n10391 , n10392 );
and ( n10394 , n10393 , n2422 );
and ( n10395 , n4231 , n2428 );
or ( n10396 , n10394 , n10395 );
buf ( n10397 , n10396 );
buf ( n10398 , n2424 );
buf ( n10399 , n2281 );
buf ( n10400 , n2280 );
not ( n10401 , n3260 );
and ( n10402 , n7339 , n5249 );
and ( n10403 , n4221 , n10237 );
or ( n10404 , n10402 , n10403 );
and ( n10405 , n10404 , n5285 );
and ( n10406 , n7350 , n5249 );
and ( n10407 , n4221 , n10237 );
or ( n10408 , n10406 , n10407 );
and ( n10409 , n10408 , n6218 );
and ( n10410 , n7361 , n5249 );
and ( n10411 , n4221 , n10237 );
or ( n10412 , n10410 , n10411 );
and ( n10413 , n10412 , n6710 );
and ( n10414 , n5717 , n5249 );
and ( n10415 , n4221 , n10237 );
or ( n10416 , n10414 , n10415 );
and ( n10417 , n10416 , n6717 );
and ( n10418 , n7373 , n5249 );
and ( n10419 , n4221 , n10237 );
or ( n10420 , n10418 , n10419 );
and ( n10421 , n10420 , n6724 );
and ( n10422 , n4221 , n9115 );
or ( n10423 , n10405 , n10409 , n10413 , n10417 , n10421 , n10422 );
and ( n10424 , n10401 , n10423 );
and ( n10425 , n4221 , n3260 );
or ( n10426 , n10424 , n10425 );
and ( n10427 , n10426 , n2422 );
and ( n10428 , n4221 , n2428 );
or ( n10429 , n10427 , n10428 );
buf ( n10430 , n10429 );
buf ( n10431 , n2424 );
buf ( n10432 , n2281 );
buf ( n10433 , n2280 );
not ( n10434 , n3260 );
and ( n10435 , n7413 , n5249 );
and ( n10436 , n4211 , n10237 );
or ( n10437 , n10435 , n10436 );
and ( n10438 , n10437 , n5285 );
and ( n10439 , n7424 , n5249 );
and ( n10440 , n4211 , n10237 );
or ( n10441 , n10439 , n10440 );
and ( n10442 , n10441 , n6218 );
and ( n10443 , n7435 , n5249 );
and ( n10444 , n4211 , n10237 );
or ( n10445 , n10443 , n10444 );
and ( n10446 , n10445 , n6710 );
and ( n10447 , n5707 , n5249 );
and ( n10448 , n4211 , n10237 );
or ( n10449 , n10447 , n10448 );
and ( n10450 , n10449 , n6717 );
and ( n10451 , n7447 , n5249 );
and ( n10452 , n4211 , n10237 );
or ( n10453 , n10451 , n10452 );
and ( n10454 , n10453 , n6724 );
and ( n10455 , n4211 , n9115 );
or ( n10456 , n10438 , n10442 , n10446 , n10450 , n10454 , n10455 );
and ( n10457 , n10434 , n10456 );
and ( n10458 , n4211 , n3260 );
or ( n10459 , n10457 , n10458 );
and ( n10460 , n10459 , n2422 );
and ( n10461 , n4211 , n2428 );
or ( n10462 , n10460 , n10461 );
buf ( n10463 , n10462 );
buf ( n10464 , n2424 );
buf ( n10465 , n2281 );
buf ( n10466 , n2280 );
not ( n10467 , n3260 );
and ( n10468 , n7487 , n5249 );
and ( n10469 , n4201 , n10237 );
or ( n10470 , n10468 , n10469 );
and ( n10471 , n10470 , n5285 );
and ( n10472 , n7498 , n5249 );
and ( n10473 , n4201 , n10237 );
or ( n10474 , n10472 , n10473 );
and ( n10475 , n10474 , n6218 );
and ( n10476 , n7509 , n5249 );
and ( n10477 , n4201 , n10237 );
or ( n10478 , n10476 , n10477 );
and ( n10479 , n10478 , n6710 );
and ( n10480 , n5697 , n5249 );
and ( n10481 , n4201 , n10237 );
or ( n10482 , n10480 , n10481 );
and ( n10483 , n10482 , n6717 );
and ( n10484 , n7521 , n5249 );
and ( n10485 , n4201 , n10237 );
or ( n10486 , n10484 , n10485 );
and ( n10487 , n10486 , n6724 );
and ( n10488 , n4201 , n9115 );
or ( n10489 , n10471 , n10475 , n10479 , n10483 , n10487 , n10488 );
and ( n10490 , n10467 , n10489 );
and ( n10491 , n4201 , n3260 );
or ( n10492 , n10490 , n10491 );
and ( n10493 , n10492 , n2422 );
and ( n10494 , n4201 , n2428 );
or ( n10495 , n10493 , n10494 );
buf ( n10496 , n10495 );
buf ( n10497 , n2424 );
buf ( n10498 , n2281 );
buf ( n10499 , n2280 );
not ( n10500 , n3260 );
and ( n10501 , n7561 , n5249 );
and ( n10502 , n4191 , n10237 );
or ( n10503 , n10501 , n10502 );
and ( n10504 , n10503 , n5285 );
and ( n10505 , n7572 , n5249 );
and ( n10506 , n4191 , n10237 );
or ( n10507 , n10505 , n10506 );
and ( n10508 , n10507 , n6218 );
and ( n10509 , n7583 , n5249 );
and ( n10510 , n4191 , n10237 );
or ( n10511 , n10509 , n10510 );
and ( n10512 , n10511 , n6710 );
and ( n10513 , n5687 , n5249 );
and ( n10514 , n4191 , n10237 );
or ( n10515 , n10513 , n10514 );
and ( n10516 , n10515 , n6717 );
and ( n10517 , n7595 , n5249 );
and ( n10518 , n4191 , n10237 );
or ( n10519 , n10517 , n10518 );
and ( n10520 , n10519 , n6724 );
and ( n10521 , n4191 , n9115 );
or ( n10522 , n10504 , n10508 , n10512 , n10516 , n10520 , n10521 );
and ( n10523 , n10500 , n10522 );
and ( n10524 , n4191 , n3260 );
or ( n10525 , n10523 , n10524 );
and ( n10526 , n10525 , n2422 );
and ( n10527 , n4191 , n2428 );
or ( n10528 , n10526 , n10527 );
buf ( n10529 , n10528 );
buf ( n10530 , n2424 );
buf ( n10531 , n2281 );
buf ( n10532 , n2280 );
not ( n10533 , n3260 );
and ( n10534 , n7635 , n5249 );
and ( n10535 , n4181 , n10237 );
or ( n10536 , n10534 , n10535 );
and ( n10537 , n10536 , n5285 );
and ( n10538 , n7646 , n5249 );
and ( n10539 , n4181 , n10237 );
or ( n10540 , n10538 , n10539 );
and ( n10541 , n10540 , n6218 );
and ( n10542 , n7657 , n5249 );
and ( n10543 , n4181 , n10237 );
or ( n10544 , n10542 , n10543 );
and ( n10545 , n10544 , n6710 );
and ( n10546 , n5677 , n5249 );
and ( n10547 , n4181 , n10237 );
or ( n10548 , n10546 , n10547 );
and ( n10549 , n10548 , n6717 );
and ( n10550 , n7669 , n5249 );
and ( n10551 , n4181 , n10237 );
or ( n10552 , n10550 , n10551 );
and ( n10553 , n10552 , n6724 );
and ( n10554 , n4181 , n9115 );
or ( n10555 , n10537 , n10541 , n10545 , n10549 , n10553 , n10554 );
and ( n10556 , n10533 , n10555 );
and ( n10557 , n4181 , n3260 );
or ( n10558 , n10556 , n10557 );
and ( n10559 , n10558 , n2422 );
and ( n10560 , n4181 , n2428 );
or ( n10561 , n10559 , n10560 );
buf ( n10562 , n10561 );
buf ( n10563 , n2424 );
buf ( n10564 , n2281 );
buf ( n10565 , n2280 );
not ( n10566 , n3260 );
and ( n10567 , n7709 , n5249 );
and ( n10568 , n4171 , n10237 );
or ( n10569 , n10567 , n10568 );
and ( n10570 , n10569 , n5285 );
and ( n10571 , n7720 , n5249 );
and ( n10572 , n4171 , n10237 );
or ( n10573 , n10571 , n10572 );
and ( n10574 , n10573 , n6218 );
and ( n10575 , n7731 , n5249 );
and ( n10576 , n4171 , n10237 );
or ( n10577 , n10575 , n10576 );
and ( n10578 , n10577 , n6710 );
and ( n10579 , n5667 , n5249 );
and ( n10580 , n4171 , n10237 );
or ( n10581 , n10579 , n10580 );
and ( n10582 , n10581 , n6717 );
and ( n10583 , n7743 , n5249 );
and ( n10584 , n4171 , n10237 );
or ( n10585 , n10583 , n10584 );
and ( n10586 , n10585 , n6724 );
and ( n10587 , n4171 , n9115 );
or ( n10588 , n10570 , n10574 , n10578 , n10582 , n10586 , n10587 );
and ( n10589 , n10566 , n10588 );
and ( n10590 , n4171 , n3260 );
or ( n10591 , n10589 , n10590 );
and ( n10592 , n10591 , n2422 );
and ( n10593 , n4171 , n2428 );
or ( n10594 , n10592 , n10593 );
buf ( n10595 , n10594 );
buf ( n10596 , n2424 );
buf ( n10597 , n2281 );
buf ( n10598 , n2280 );
not ( n10599 , n3260 );
and ( n10600 , n7783 , n5249 );
and ( n10601 , n4161 , n10237 );
or ( n10602 , n10600 , n10601 );
and ( n10603 , n10602 , n5285 );
and ( n10604 , n7794 , n5249 );
and ( n10605 , n4161 , n10237 );
or ( n10606 , n10604 , n10605 );
and ( n10607 , n10606 , n6218 );
and ( n10608 , n7805 , n5249 );
and ( n10609 , n4161 , n10237 );
or ( n10610 , n10608 , n10609 );
and ( n10611 , n10610 , n6710 );
and ( n10612 , n5657 , n5249 );
and ( n10613 , n4161 , n10237 );
or ( n10614 , n10612 , n10613 );
and ( n10615 , n10614 , n6717 );
and ( n10616 , n7817 , n5249 );
and ( n10617 , n4161 , n10237 );
or ( n10618 , n10616 , n10617 );
and ( n10619 , n10618 , n6724 );
and ( n10620 , n4161 , n9115 );
or ( n10621 , n10603 , n10607 , n10611 , n10615 , n10619 , n10620 );
and ( n10622 , n10599 , n10621 );
and ( n10623 , n4161 , n3260 );
or ( n10624 , n10622 , n10623 );
and ( n10625 , n10624 , n2422 );
and ( n10626 , n4161 , n2428 );
or ( n10627 , n10625 , n10626 );
buf ( n10628 , n10627 );
buf ( n10629 , n2424 );
buf ( n10630 , n2281 );
buf ( n10631 , n2280 );
not ( n10632 , n3260 );
and ( n10633 , n7857 , n5249 );
and ( n10634 , n4151 , n10237 );
or ( n10635 , n10633 , n10634 );
and ( n10636 , n10635 , n5285 );
and ( n10637 , n7868 , n5249 );
and ( n10638 , n4151 , n10237 );
or ( n10639 , n10637 , n10638 );
and ( n10640 , n10639 , n6218 );
and ( n10641 , n7879 , n5249 );
and ( n10642 , n4151 , n10237 );
or ( n10643 , n10641 , n10642 );
and ( n10644 , n10643 , n6710 );
and ( n10645 , n5647 , n5249 );
and ( n10646 , n4151 , n10237 );
or ( n10647 , n10645 , n10646 );
and ( n10648 , n10647 , n6717 );
and ( n10649 , n7891 , n5249 );
and ( n10650 , n4151 , n10237 );
or ( n10651 , n10649 , n10650 );
and ( n10652 , n10651 , n6724 );
and ( n10653 , n4151 , n9115 );
or ( n10654 , n10636 , n10640 , n10644 , n10648 , n10652 , n10653 );
and ( n10655 , n10632 , n10654 );
and ( n10656 , n4151 , n3260 );
or ( n10657 , n10655 , n10656 );
and ( n10658 , n10657 , n2422 );
and ( n10659 , n4151 , n2428 );
or ( n10660 , n10658 , n10659 );
buf ( n10661 , n10660 );
buf ( n10662 , n2424 );
buf ( n10663 , n2281 );
buf ( n10664 , n2280 );
not ( n10665 , n3260 );
and ( n10666 , n7931 , n5249 );
and ( n10667 , n4141 , n10237 );
or ( n10668 , n10666 , n10667 );
and ( n10669 , n10668 , n5285 );
and ( n10670 , n7942 , n5249 );
and ( n10671 , n4141 , n10237 );
or ( n10672 , n10670 , n10671 );
and ( n10673 , n10672 , n6218 );
and ( n10674 , n7953 , n5249 );
and ( n10675 , n4141 , n10237 );
or ( n10676 , n10674 , n10675 );
and ( n10677 , n10676 , n6710 );
and ( n10678 , n5637 , n5249 );
and ( n10679 , n4141 , n10237 );
or ( n10680 , n10678 , n10679 );
and ( n10681 , n10680 , n6717 );
and ( n10682 , n7965 , n5249 );
and ( n10683 , n4141 , n10237 );
or ( n10684 , n10682 , n10683 );
and ( n10685 , n10684 , n6724 );
and ( n10686 , n4141 , n9115 );
or ( n10687 , n10669 , n10673 , n10677 , n10681 , n10685 , n10686 );
and ( n10688 , n10665 , n10687 );
and ( n10689 , n4141 , n3260 );
or ( n10690 , n10688 , n10689 );
and ( n10691 , n10690 , n2422 );
and ( n10692 , n4141 , n2428 );
or ( n10693 , n10691 , n10692 );
buf ( n10694 , n10693 );
buf ( n10695 , n2424 );
buf ( n10696 , n2281 );
buf ( n10697 , n2280 );
not ( n10698 , n3260 );
and ( n10699 , n8005 , n5249 );
and ( n10700 , n4131 , n10237 );
or ( n10701 , n10699 , n10700 );
and ( n10702 , n10701 , n5285 );
and ( n10703 , n8016 , n5249 );
and ( n10704 , n4131 , n10237 );
or ( n10705 , n10703 , n10704 );
and ( n10706 , n10705 , n6218 );
and ( n10707 , n8027 , n5249 );
and ( n10708 , n4131 , n10237 );
or ( n10709 , n10707 , n10708 );
and ( n10710 , n10709 , n6710 );
and ( n10711 , n5627 , n5249 );
and ( n10712 , n4131 , n10237 );
or ( n10713 , n10711 , n10712 );
and ( n10714 , n10713 , n6717 );
and ( n10715 , n8039 , n5249 );
and ( n10716 , n4131 , n10237 );
or ( n10717 , n10715 , n10716 );
and ( n10718 , n10717 , n6724 );
and ( n10719 , n4131 , n9115 );
or ( n10720 , n10702 , n10706 , n10710 , n10714 , n10718 , n10719 );
and ( n10721 , n10698 , n10720 );
and ( n10722 , n4131 , n3260 );
or ( n10723 , n10721 , n10722 );
and ( n10724 , n10723 , n2422 );
and ( n10725 , n4131 , n2428 );
or ( n10726 , n10724 , n10725 );
buf ( n10727 , n10726 );
buf ( n10728 , n2424 );
buf ( n10729 , n2281 );
buf ( n10730 , n2280 );
not ( n10731 , n3260 );
and ( n10732 , n8079 , n5249 );
and ( n10733 , n4121 , n10237 );
or ( n10734 , n10732 , n10733 );
and ( n10735 , n10734 , n5285 );
and ( n10736 , n8090 , n5249 );
and ( n10737 , n4121 , n10237 );
or ( n10738 , n10736 , n10737 );
and ( n10739 , n10738 , n6218 );
and ( n10740 , n8101 , n5249 );
and ( n10741 , n4121 , n10237 );
or ( n10742 , n10740 , n10741 );
and ( n10743 , n10742 , n6710 );
and ( n10744 , n5617 , n5249 );
and ( n10745 , n4121 , n10237 );
or ( n10746 , n10744 , n10745 );
and ( n10747 , n10746 , n6717 );
and ( n10748 , n8113 , n5249 );
and ( n10749 , n4121 , n10237 );
or ( n10750 , n10748 , n10749 );
and ( n10751 , n10750 , n6724 );
and ( n10752 , n4121 , n9115 );
or ( n10753 , n10735 , n10739 , n10743 , n10747 , n10751 , n10752 );
and ( n10754 , n10731 , n10753 );
and ( n10755 , n4121 , n3260 );
or ( n10756 , n10754 , n10755 );
and ( n10757 , n10756 , n2422 );
and ( n10758 , n4121 , n2428 );
or ( n10759 , n10757 , n10758 );
buf ( n10760 , n10759 );
buf ( n10761 , n2424 );
buf ( n10762 , n2281 );
buf ( n10763 , n2280 );
not ( n10764 , n3260 );
and ( n10765 , n8153 , n5249 );
and ( n10766 , n4111 , n10237 );
or ( n10767 , n10765 , n10766 );
and ( n10768 , n10767 , n5285 );
and ( n10769 , n8164 , n5249 );
and ( n10770 , n4111 , n10237 );
or ( n10771 , n10769 , n10770 );
and ( n10772 , n10771 , n6218 );
and ( n10773 , n8175 , n5249 );
and ( n10774 , n4111 , n10237 );
or ( n10775 , n10773 , n10774 );
and ( n10776 , n10775 , n6710 );
and ( n10777 , n5607 , n5249 );
and ( n10778 , n4111 , n10237 );
or ( n10779 , n10777 , n10778 );
and ( n10780 , n10779 , n6717 );
and ( n10781 , n8187 , n5249 );
and ( n10782 , n4111 , n10237 );
or ( n10783 , n10781 , n10782 );
and ( n10784 , n10783 , n6724 );
and ( n10785 , n4111 , n9115 );
or ( n10786 , n10768 , n10772 , n10776 , n10780 , n10784 , n10785 );
and ( n10787 , n10764 , n10786 );
and ( n10788 , n4111 , n3260 );
or ( n10789 , n10787 , n10788 );
and ( n10790 , n10789 , n2422 );
and ( n10791 , n4111 , n2428 );
or ( n10792 , n10790 , n10791 );
buf ( n10793 , n10792 );
buf ( n10794 , n2424 );
buf ( n10795 , n2281 );
buf ( n10796 , n2280 );
not ( n10797 , n3260 );
and ( n10798 , n8227 , n5249 );
and ( n10799 , n4101 , n10237 );
or ( n10800 , n10798 , n10799 );
and ( n10801 , n10800 , n5285 );
and ( n10802 , n8238 , n5249 );
and ( n10803 , n4101 , n10237 );
or ( n10804 , n10802 , n10803 );
and ( n10805 , n10804 , n6218 );
and ( n10806 , n8249 , n5249 );
and ( n10807 , n4101 , n10237 );
or ( n10808 , n10806 , n10807 );
and ( n10809 , n10808 , n6710 );
and ( n10810 , n5597 , n5249 );
and ( n10811 , n4101 , n10237 );
or ( n10812 , n10810 , n10811 );
and ( n10813 , n10812 , n6717 );
and ( n10814 , n8261 , n5249 );
and ( n10815 , n4101 , n10237 );
or ( n10816 , n10814 , n10815 );
and ( n10817 , n10816 , n6724 );
and ( n10818 , n4101 , n9115 );
or ( n10819 , n10801 , n10805 , n10809 , n10813 , n10817 , n10818 );
and ( n10820 , n10797 , n10819 );
and ( n10821 , n4101 , n3260 );
or ( n10822 , n10820 , n10821 );
and ( n10823 , n10822 , n2422 );
and ( n10824 , n4101 , n2428 );
or ( n10825 , n10823 , n10824 );
buf ( n10826 , n10825 );
buf ( n10827 , n2424 );
buf ( n10828 , n2281 );
buf ( n10829 , n2280 );
not ( n10830 , n3260 );
and ( n10831 , n8301 , n5249 );
and ( n10832 , n4091 , n10237 );
or ( n10833 , n10831 , n10832 );
and ( n10834 , n10833 , n5285 );
and ( n10835 , n8312 , n5249 );
and ( n10836 , n4091 , n10237 );
or ( n10837 , n10835 , n10836 );
and ( n10838 , n10837 , n6218 );
and ( n10839 , n8323 , n5249 );
and ( n10840 , n4091 , n10237 );
or ( n10841 , n10839 , n10840 );
and ( n10842 , n10841 , n6710 );
and ( n10843 , n5587 , n5249 );
and ( n10844 , n4091 , n10237 );
or ( n10845 , n10843 , n10844 );
and ( n10846 , n10845 , n6717 );
and ( n10847 , n8335 , n5249 );
and ( n10848 , n4091 , n10237 );
or ( n10849 , n10847 , n10848 );
and ( n10850 , n10849 , n6724 );
and ( n10851 , n4091 , n9115 );
or ( n10852 , n10834 , n10838 , n10842 , n10846 , n10850 , n10851 );
and ( n10853 , n10830 , n10852 );
and ( n10854 , n4091 , n3260 );
or ( n10855 , n10853 , n10854 );
and ( n10856 , n10855 , n2422 );
and ( n10857 , n4091 , n2428 );
or ( n10858 , n10856 , n10857 );
buf ( n10859 , n10858 );
buf ( n10860 , n2424 );
buf ( n10861 , n2281 );
buf ( n10862 , n2280 );
not ( n10863 , n3260 );
and ( n10864 , n8375 , n5249 );
and ( n10865 , n4081 , n10237 );
or ( n10866 , n10864 , n10865 );
and ( n10867 , n10866 , n5285 );
and ( n10868 , n8386 , n5249 );
and ( n10869 , n4081 , n10237 );
or ( n10870 , n10868 , n10869 );
and ( n10871 , n10870 , n6218 );
and ( n10872 , n8397 , n5249 );
and ( n10873 , n4081 , n10237 );
or ( n10874 , n10872 , n10873 );
and ( n10875 , n10874 , n6710 );
and ( n10876 , n5577 , n5249 );
and ( n10877 , n4081 , n10237 );
or ( n10878 , n10876 , n10877 );
and ( n10879 , n10878 , n6717 );
and ( n10880 , n8409 , n5249 );
and ( n10881 , n4081 , n10237 );
or ( n10882 , n10880 , n10881 );
and ( n10883 , n10882 , n6724 );
and ( n10884 , n4081 , n9115 );
or ( n10885 , n10867 , n10871 , n10875 , n10879 , n10883 , n10884 );
and ( n10886 , n10863 , n10885 );
and ( n10887 , n4081 , n3260 );
or ( n10888 , n10886 , n10887 );
and ( n10889 , n10888 , n2422 );
and ( n10890 , n4081 , n2428 );
or ( n10891 , n10889 , n10890 );
buf ( n10892 , n10891 );
buf ( n10893 , n2424 );
buf ( n10894 , n2281 );
buf ( n10895 , n2280 );
not ( n10896 , n3260 );
and ( n10897 , n8449 , n5249 );
and ( n10898 , n4071 , n10237 );
or ( n10899 , n10897 , n10898 );
and ( n10900 , n10899 , n5285 );
and ( n10901 , n8460 , n5249 );
and ( n10902 , n4071 , n10237 );
or ( n10903 , n10901 , n10902 );
and ( n10904 , n10903 , n6218 );
and ( n10905 , n8471 , n5249 );
and ( n10906 , n4071 , n10237 );
or ( n10907 , n10905 , n10906 );
and ( n10908 , n10907 , n6710 );
and ( n10909 , n5529 , n5249 );
and ( n10910 , n4071 , n10237 );
or ( n10911 , n10909 , n10910 );
and ( n10912 , n10911 , n6717 );
and ( n10913 , n8483 , n5249 );
and ( n10914 , n4071 , n10237 );
or ( n10915 , n10913 , n10914 );
and ( n10916 , n10915 , n6724 );
and ( n10917 , n4071 , n9115 );
or ( n10918 , n10900 , n10904 , n10908 , n10912 , n10916 , n10917 );
and ( n10919 , n10896 , n10918 );
and ( n10920 , n4071 , n3260 );
or ( n10921 , n10919 , n10920 );
and ( n10922 , n10921 , n2422 );
and ( n10923 , n4071 , n2428 );
or ( n10924 , n10922 , n10923 );
buf ( n10925 , n10924 );
buf ( n10926 , n2424 );
buf ( n10927 , n2281 );
buf ( n10928 , n2280 );
not ( n10929 , n3260 );
and ( n10930 , n8523 , n5249 );
and ( n10931 , n4061 , n10237 );
or ( n10932 , n10930 , n10931 );
and ( n10933 , n10932 , n5285 );
and ( n10934 , n8534 , n5249 );
and ( n10935 , n4061 , n10237 );
or ( n10936 , n10934 , n10935 );
and ( n10937 , n10936 , n6218 );
and ( n10938 , n8545 , n5249 );
and ( n10939 , n4061 , n10237 );
or ( n10940 , n10938 , n10939 );
and ( n10941 , n10940 , n6710 );
and ( n10942 , n5526 , n5249 );
and ( n10943 , n4061 , n10237 );
or ( n10944 , n10942 , n10943 );
and ( n10945 , n10944 , n6717 );
and ( n10946 , n8557 , n5249 );
and ( n10947 , n4061 , n10237 );
or ( n10948 , n10946 , n10947 );
and ( n10949 , n10948 , n6724 );
and ( n10950 , n4061 , n9115 );
or ( n10951 , n10933 , n10937 , n10941 , n10945 , n10949 , n10950 );
and ( n10952 , n10929 , n10951 );
and ( n10953 , n4061 , n3260 );
or ( n10954 , n10952 , n10953 );
and ( n10955 , n10954 , n2422 );
and ( n10956 , n4061 , n2428 );
or ( n10957 , n10955 , n10956 );
buf ( n10958 , n10957 );
buf ( n10959 , n2424 );
buf ( n10960 , n2281 );
buf ( n10961 , n2280 );
not ( n10962 , n3260 );
and ( n10963 , n8597 , n5249 );
and ( n10964 , n4051 , n10237 );
or ( n10965 , n10963 , n10964 );
and ( n10966 , n10965 , n5285 );
and ( n10967 , n8608 , n5249 );
and ( n10968 , n4051 , n10237 );
or ( n10969 , n10967 , n10968 );
and ( n10970 , n10969 , n6218 );
and ( n10971 , n8619 , n5249 );
and ( n10972 , n4051 , n10237 );
or ( n10973 , n10971 , n10972 );
and ( n10974 , n10973 , n6710 );
and ( n10975 , n5523 , n5249 );
and ( n10976 , n4051 , n10237 );
or ( n10977 , n10975 , n10976 );
and ( n10978 , n10977 , n6717 );
and ( n10979 , n8631 , n5249 );
and ( n10980 , n4051 , n10237 );
or ( n10981 , n10979 , n10980 );
and ( n10982 , n10981 , n6724 );
and ( n10983 , n4051 , n9115 );
or ( n10984 , n10966 , n10970 , n10974 , n10978 , n10982 , n10983 );
and ( n10985 , n10962 , n10984 );
and ( n10986 , n4051 , n3260 );
or ( n10987 , n10985 , n10986 );
and ( n10988 , n10987 , n2422 );
and ( n10989 , n4051 , n2428 );
or ( n10990 , n10988 , n10989 );
buf ( n10991 , n10990 );
buf ( n10992 , n2424 );
buf ( n10993 , n2281 );
buf ( n10994 , n2280 );
not ( n10995 , n3260 );
and ( n10996 , n8671 , n5249 );
and ( n10997 , n4041 , n10237 );
or ( n10998 , n10996 , n10997 );
and ( n10999 , n10998 , n5285 );
and ( n11000 , n8682 , n5249 );
and ( n11001 , n4041 , n10237 );
or ( n11002 , n11000 , n11001 );
and ( n11003 , n11002 , n6218 );
and ( n11004 , n8693 , n5249 );
and ( n11005 , n4041 , n10237 );
or ( n11006 , n11004 , n11005 );
and ( n11007 , n11006 , n6710 );
and ( n11008 , n5520 , n5249 );
and ( n11009 , n4041 , n10237 );
or ( n11010 , n11008 , n11009 );
and ( n11011 , n11010 , n6717 );
and ( n11012 , n8705 , n5249 );
and ( n11013 , n4041 , n10237 );
or ( n11014 , n11012 , n11013 );
and ( n11015 , n11014 , n6724 );
and ( n11016 , n4041 , n9115 );
or ( n11017 , n10999 , n11003 , n11007 , n11011 , n11015 , n11016 );
and ( n11018 , n10995 , n11017 );
and ( n11019 , n4041 , n3260 );
or ( n11020 , n11018 , n11019 );
and ( n11021 , n11020 , n2422 );
and ( n11022 , n4041 , n2428 );
or ( n11023 , n11021 , n11022 );
buf ( n11024 , n11023 );
buf ( n11025 , n2424 );
buf ( n11026 , n2281 );
buf ( n11027 , n2280 );
not ( n11028 , n3260 );
and ( n11029 , n8745 , n5249 );
and ( n11030 , n4031 , n10237 );
or ( n11031 , n11029 , n11030 );
and ( n11032 , n11031 , n5285 );
and ( n11033 , n8756 , n5249 );
and ( n11034 , n4031 , n10237 );
or ( n11035 , n11033 , n11034 );
and ( n11036 , n11035 , n6218 );
and ( n11037 , n8767 , n5249 );
and ( n11038 , n4031 , n10237 );
or ( n11039 , n11037 , n11038 );
and ( n11040 , n11039 , n6710 );
and ( n11041 , n5517 , n5249 );
and ( n11042 , n4031 , n10237 );
or ( n11043 , n11041 , n11042 );
and ( n11044 , n11043 , n6717 );
and ( n11045 , n8779 , n5249 );
and ( n11046 , n4031 , n10237 );
or ( n11047 , n11045 , n11046 );
and ( n11048 , n11047 , n6724 );
and ( n11049 , n4031 , n9115 );
or ( n11050 , n11032 , n11036 , n11040 , n11044 , n11048 , n11049 );
and ( n11051 , n11028 , n11050 );
and ( n11052 , n4031 , n3260 );
or ( n11053 , n11051 , n11052 );
and ( n11054 , n11053 , n2422 );
and ( n11055 , n4031 , n2428 );
or ( n11056 , n11054 , n11055 );
buf ( n11057 , n11056 );
buf ( n11058 , n2424 );
buf ( n11059 , n2281 );
buf ( n11060 , n2280 );
not ( n11061 , n3260 );
and ( n11062 , n8819 , n5249 );
and ( n11063 , n4021 , n10237 );
or ( n11064 , n11062 , n11063 );
and ( n11065 , n11064 , n5285 );
and ( n11066 , n8830 , n5249 );
and ( n11067 , n4021 , n10237 );
or ( n11068 , n11066 , n11067 );
and ( n11069 , n11068 , n6218 );
and ( n11070 , n8841 , n5249 );
and ( n11071 , n4021 , n10237 );
or ( n11072 , n11070 , n11071 );
and ( n11073 , n11072 , n6710 );
and ( n11074 , n5514 , n5249 );
and ( n11075 , n4021 , n10237 );
or ( n11076 , n11074 , n11075 );
and ( n11077 , n11076 , n6717 );
and ( n11078 , n8853 , n5249 );
and ( n11079 , n4021 , n10237 );
or ( n11080 , n11078 , n11079 );
and ( n11081 , n11080 , n6724 );
and ( n11082 , n4021 , n9115 );
or ( n11083 , n11065 , n11069 , n11073 , n11077 , n11081 , n11082 );
and ( n11084 , n11061 , n11083 );
and ( n11085 , n4021 , n3260 );
or ( n11086 , n11084 , n11085 );
and ( n11087 , n11086 , n2422 );
and ( n11088 , n4021 , n2428 );
or ( n11089 , n11087 , n11088 );
buf ( n11090 , n11089 );
buf ( n11091 , n2424 );
buf ( n11092 , n2281 );
buf ( n11093 , n2280 );
not ( n11094 , n3260 );
and ( n11095 , n8893 , n5249 );
and ( n11096 , n4011 , n10237 );
or ( n11097 , n11095 , n11096 );
and ( n11098 , n11097 , n5285 );
and ( n11099 , n8904 , n5249 );
and ( n11100 , n4011 , n10237 );
or ( n11101 , n11099 , n11100 );
and ( n11102 , n11101 , n6218 );
and ( n11103 , n8915 , n5249 );
and ( n11104 , n4011 , n10237 );
or ( n11105 , n11103 , n11104 );
and ( n11106 , n11105 , n6710 );
and ( n11107 , n5511 , n5249 );
and ( n11108 , n4011 , n10237 );
or ( n11109 , n11107 , n11108 );
and ( n11110 , n11109 , n6717 );
and ( n11111 , n8927 , n5249 );
and ( n11112 , n4011 , n10237 );
or ( n11113 , n11111 , n11112 );
and ( n11114 , n11113 , n6724 );
and ( n11115 , n4011 , n9115 );
or ( n11116 , n11098 , n11102 , n11106 , n11110 , n11114 , n11115 );
and ( n11117 , n11094 , n11116 );
and ( n11118 , n4011 , n3260 );
or ( n11119 , n11117 , n11118 );
and ( n11120 , n11119 , n2422 );
and ( n11121 , n4011 , n2428 );
or ( n11122 , n11120 , n11121 );
buf ( n11123 , n11122 );
buf ( n11124 , n2424 );
buf ( n11125 , n2281 );
buf ( n11126 , n2280 );
not ( n11127 , n3260 );
and ( n11128 , n8967 , n5249 );
and ( n11129 , n4001 , n10237 );
or ( n11130 , n11128 , n11129 );
and ( n11131 , n11130 , n5285 );
and ( n11132 , n8978 , n5249 );
and ( n11133 , n4001 , n10237 );
or ( n11134 , n11132 , n11133 );
and ( n11135 , n11134 , n6218 );
and ( n11136 , n8989 , n5249 );
and ( n11137 , n4001 , n10237 );
or ( n11138 , n11136 , n11137 );
and ( n11139 , n11138 , n6710 );
and ( n11140 , n5508 , n5249 );
and ( n11141 , n4001 , n10237 );
or ( n11142 , n11140 , n11141 );
and ( n11143 , n11142 , n6717 );
and ( n11144 , n9001 , n5249 );
and ( n11145 , n4001 , n10237 );
or ( n11146 , n11144 , n11145 );
and ( n11147 , n11146 , n6724 );
and ( n11148 , n4001 , n9115 );
or ( n11149 , n11131 , n11135 , n11139 , n11143 , n11147 , n11148 );
and ( n11150 , n11127 , n11149 );
and ( n11151 , n4001 , n3260 );
or ( n11152 , n11150 , n11151 );
and ( n11153 , n11152 , n2422 );
and ( n11154 , n4001 , n2428 );
or ( n11155 , n11153 , n11154 );
buf ( n11156 , n11155 );
buf ( n11157 , n2424 );
buf ( n11158 , n2281 );
buf ( n11159 , n2280 );
not ( n11160 , n3260 );
and ( n11161 , n9041 , n5249 );
and ( n11162 , n3991 , n10237 );
or ( n11163 , n11161 , n11162 );
and ( n11164 , n11163 , n5285 );
and ( n11165 , n9052 , n5249 );
and ( n11166 , n3991 , n10237 );
or ( n11167 , n11165 , n11166 );
and ( n11168 , n11167 , n6218 );
and ( n11169 , n9063 , n5249 );
and ( n11170 , n3991 , n10237 );
or ( n11171 , n11169 , n11170 );
and ( n11172 , n11171 , n6710 );
and ( n11173 , n5505 , n5249 );
and ( n11174 , n3991 , n10237 );
or ( n11175 , n11173 , n11174 );
and ( n11176 , n11175 , n6717 );
and ( n11177 , n9075 , n5249 );
and ( n11178 , n3991 , n10237 );
or ( n11179 , n11177 , n11178 );
and ( n11180 , n11179 , n6724 );
and ( n11181 , n3991 , n9115 );
or ( n11182 , n11164 , n11168 , n11172 , n11176 , n11180 , n11181 );
and ( n11183 , n11160 , n11182 );
and ( n11184 , n3991 , n3260 );
or ( n11185 , n11183 , n11184 );
and ( n11186 , n11185 , n2422 );
nand ( n11187 , n3991 , n2428 );
or ( n11188 , n11186 , n11187 );
buf ( n11189 , n11188 );
buf ( n11190 , n2424 );
buf ( n11191 , n2281 );
buf ( n11192 , n2280 );
not ( n11193 , n3260 );
and ( n11194 , n10078 , n5249 );
and ( n11195 , n3981 , n10237 );
or ( n11196 , n11194 , n11195 );
and ( n11197 , n11196 , n5285 );
and ( n11198 , n10089 , n5249 );
and ( n11199 , n3981 , n10237 );
or ( n11200 , n11198 , n11199 );
and ( n11201 , n11200 , n6218 );
and ( n11202 , n10100 , n5249 );
and ( n11203 , n3981 , n10237 );
or ( n11204 , n11202 , n11203 );
and ( n11205 , n11204 , n6710 );
and ( n11206 , n5502 , n5249 );
and ( n11207 , n3981 , n10237 );
or ( n11208 , n11206 , n11207 );
and ( n11209 , n11208 , n6717 );
and ( n11210 , n10111 , n5249 );
and ( n11211 , n3981 , n10237 );
or ( n11212 , n11210 , n11211 );
and ( n11213 , n11212 , n6724 );
and ( n11214 , n3981 , n9115 );
or ( n11215 , n11197 , n11201 , n11205 , n11209 , n11213 , n11214 );
and ( n11216 , n11193 , n11215 );
and ( n11217 , n3981 , n3260 );
or ( n11218 , n11216 , n11217 );
and ( n11219 , n11218 , n2422 );
and ( n11220 , n3981 , n2428 );
or ( n11221 , n11219 , n11220 );
buf ( n11222 , n11221 );
buf ( n11223 , n2424 );
buf ( n11224 , n2281 );
buf ( n11225 , n2280 );
not ( n11226 , n3260 );
and ( n11227 , n10147 , n5249 );
and ( n11228 , n3817 , n10237 );
or ( n11229 , n11227 , n11228 );
and ( n11230 , n11229 , n5285 );
and ( n11231 , n10156 , n5249 );
and ( n11232 , n3817 , n10237 );
or ( n11233 , n11231 , n11232 );
and ( n11234 , n11233 , n6218 );
and ( n11235 , n10165 , n5249 );
and ( n11236 , n3817 , n10237 );
or ( n11237 , n11235 , n11236 );
and ( n11238 , n11237 , n6710 );
and ( n11239 , n5499 , n5249 );
and ( n11240 , n3817 , n10237 );
or ( n11241 , n11239 , n11240 );
and ( n11242 , n11241 , n6717 );
and ( n11243 , n10176 , n5249 );
and ( n11244 , n3817 , n10237 );
or ( n11245 , n11243 , n11244 );
and ( n11246 , n11245 , n6724 );
and ( n11247 , n3817 , n9115 );
or ( n11248 , n11230 , n11234 , n11238 , n11242 , n11246 , n11247 );
and ( n11249 , n11226 , n11248 );
and ( n11250 , n3817 , n3260 );
or ( n11251 , n11249 , n11250 );
and ( n11252 , n11251 , n2422 );
and ( n11253 , n3817 , n2428 );
or ( n11254 , n11252 , n11253 );
buf ( n11255 , n11254 );
buf ( n11256 , n2424 );
buf ( n11257 , n2281 );
buf ( n11258 , n2280 );
not ( n11259 , n3260 );
and ( n11260 , n10201 , n5249 );
and ( n11261 , n3767 , n10237 );
or ( n11262 , n11260 , n11261 );
and ( n11263 , n11262 , n5285 );
and ( n11264 , n3767 , n10237 );
and ( n11265 , n11264 , n6218 );
and ( n11266 , n3767 , n10237 );
and ( n11267 , n11266 , n6710 );
and ( n11268 , n5496 , n5249 );
and ( n11269 , n3767 , n10237 );
or ( n11270 , n11268 , n11269 );
and ( n11271 , n11270 , n6717 );
and ( n11272 , n10216 , n5249 );
and ( n11273 , n3767 , n10237 );
or ( n11274 , n11272 , n11273 );
and ( n11275 , n11274 , n6724 );
and ( n11276 , n3767 , n9115 );
or ( n11277 , n11263 , n11265 , n11267 , n11271 , n11275 , n11276 );
and ( n11278 , n11259 , n11277 );
and ( n11279 , n3767 , n3260 );
or ( n11280 , n11278 , n11279 );
and ( n11281 , n11280 , n2422 );
and ( n11282 , n3767 , n2428 );
or ( n11283 , n11281 , n11282 );
buf ( n11284 , n11283 );
buf ( n11285 , n2424 );
buf ( n11286 , n2281 );
buf ( n11287 , n2280 );
not ( n11288 , n3066 );
not ( n11289 , n3259 );
and ( n11290 , n10133 , n5289 );
or ( n11291 , n5152 , n5154 );
or ( n11292 , n11291 , n5287 );
and ( n11293 , n3290 , n11292 );
or ( n11294 , n11290 , n11293 );
and ( n11295 , n11294 , n5285 );
or ( n11296 , n6719 , n6724 );
or ( n11297 , n11296 , n6715 );
or ( n11298 , n11297 , n6716 );
or ( n11299 , n11298 , n6704 );
or ( n11300 , n11299 , n6705 );
or ( n11301 , n11300 , n6212 );
or ( n11302 , n11301 , n6213 );
or ( n11303 , n11302 , n6707 );
or ( n11304 , n11303 , n6215 );
or ( n11305 , n11304 , n6709 );
or ( n11306 , n11305 , n6217 );
or ( n11307 , n11306 , n3631 );
and ( n11308 , n3290 , n11307 );
or ( n11309 , n11295 , n11308 );
and ( n11310 , n11289 , n11309 );
and ( n11311 , n3290 , n3259 );
or ( n11312 , n11310 , n11311 );
and ( n11313 , n11288 , n11312 );
not ( n11314 , n3770 );
and ( n11315 , n11314 , n3819 );
not ( n11316 , n11315 );
and ( n11317 , n11316 , n3770 );
xnor ( n11318 , n3770 , n3819 );
and ( n11319 , n11318 , n11315 );
or ( n11320 , n11317 , n11319 );
xor ( n11321 , n11320 , n5496 );
not ( n11322 , n11321 );
not ( n11323 , n11315 );
and ( n11324 , n11323 , n3819 );
not ( n11325 , n3819 );
and ( n11326 , n11325 , n11315 );
or ( n11327 , n11324 , n11326 );
not ( n11328 , n11327 );
and ( n11329 , n11328 , n5499 );
not ( n11330 , n3983 );
and ( n11331 , n11330 , n5502 );
not ( n11332 , n3993 );
and ( n11333 , n11332 , n5505 );
not ( n11334 , n4003 );
and ( n11335 , n11334 , n5508 );
not ( n11336 , n4013 );
and ( n11337 , n11336 , n5511 );
not ( n11338 , n4023 );
and ( n11339 , n11338 , n5514 );
not ( n11340 , n4033 );
and ( n11341 , n11340 , n5517 );
not ( n11342 , n4043 );
and ( n11343 , n11342 , n5520 );
not ( n11344 , n4053 );
and ( n11345 , n11344 , n5523 );
not ( n11346 , n4063 );
and ( n11347 , n11346 , n5526 );
not ( n11348 , n4073 );
and ( n11349 , n11348 , n5529 );
not ( n11350 , n4083 );
and ( n11351 , n11350 , n5577 );
not ( n11352 , n4093 );
and ( n11353 , n11352 , n5587 );
not ( n11354 , n4103 );
and ( n11355 , n11354 , n5597 );
not ( n11356 , n4113 );
and ( n11357 , n11356 , n5607 );
not ( n11358 , n4123 );
and ( n11359 , n11358 , n5617 );
not ( n11360 , n4133 );
and ( n11361 , n11360 , n5627 );
not ( n11362 , n4143 );
and ( n11363 , n11362 , n5637 );
not ( n11364 , n4153 );
and ( n11365 , n11364 , n5647 );
not ( n11366 , n4163 );
and ( n11367 , n11366 , n5657 );
not ( n11368 , n4173 );
and ( n11369 , n11368 , n5667 );
not ( n11370 , n4183 );
and ( n11371 , n11370 , n5677 );
not ( n11372 , n4193 );
and ( n11373 , n11372 , n5687 );
not ( n11374 , n4203 );
and ( n11375 , n11374 , n5697 );
not ( n11376 , n4213 );
and ( n11377 , n11376 , n5707 );
not ( n11378 , n4223 );
and ( n11379 , n11378 , n5717 );
not ( n11380 , n4233 );
and ( n11381 , n11380 , n5727 );
not ( n11382 , n4243 );
and ( n11383 , n11382 , n5737 );
not ( n11384 , n4257 );
and ( n11385 , n11384 , n5747 );
not ( n11386 , n3785 );
and ( n11387 , n11386 , n5757 );
not ( n11388 , n3795 );
and ( n11389 , n11388 , n5492 );
xnor ( n11390 , n3785 , n5757 );
and ( n11391 , n11389 , n11390 );
or ( n11392 , n11387 , n11391 );
xnor ( n11393 , n4257 , n5747 );
and ( n11394 , n11392 , n11393 );
or ( n11395 , n11385 , n11394 );
xnor ( n11396 , n4243 , n5737 );
and ( n11397 , n11395 , n11396 );
or ( n11398 , n11383 , n11397 );
xnor ( n11399 , n4233 , n5727 );
and ( n11400 , n11398 , n11399 );
or ( n11401 , n11381 , n11400 );
xnor ( n11402 , n4223 , n5717 );
and ( n11403 , n11401 , n11402 );
or ( n11404 , n11379 , n11403 );
xnor ( n11405 , n4213 , n5707 );
and ( n11406 , n11404 , n11405 );
or ( n11407 , n11377 , n11406 );
xnor ( n11408 , n4203 , n5697 );
and ( n11409 , n11407 , n11408 );
or ( n11410 , n11375 , n11409 );
xnor ( n11411 , n4193 , n5687 );
and ( n11412 , n11410 , n11411 );
or ( n11413 , n11373 , n11412 );
xnor ( n11414 , n4183 , n5677 );
and ( n11415 , n11413 , n11414 );
or ( n11416 , n11371 , n11415 );
xnor ( n11417 , n4173 , n5667 );
and ( n11418 , n11416 , n11417 );
or ( n11419 , n11369 , n11418 );
xnor ( n11420 , n4163 , n5657 );
and ( n11421 , n11419 , n11420 );
or ( n11422 , n11367 , n11421 );
xnor ( n11423 , n4153 , n5647 );
and ( n11424 , n11422 , n11423 );
or ( n11425 , n11365 , n11424 );
xnor ( n11426 , n4143 , n5637 );
and ( n11427 , n11425 , n11426 );
or ( n11428 , n11363 , n11427 );
xnor ( n11429 , n4133 , n5627 );
and ( n11430 , n11428 , n11429 );
or ( n11431 , n11361 , n11430 );
xnor ( n11432 , n4123 , n5617 );
and ( n11433 , n11431 , n11432 );
or ( n11434 , n11359 , n11433 );
xnor ( n11435 , n4113 , n5607 );
and ( n11436 , n11434 , n11435 );
or ( n11437 , n11357 , n11436 );
xnor ( n11438 , n4103 , n5597 );
and ( n11439 , n11437 , n11438 );
or ( n11440 , n11355 , n11439 );
xnor ( n11441 , n4093 , n5587 );
and ( n11442 , n11440 , n11441 );
or ( n11443 , n11353 , n11442 );
xnor ( n11444 , n4083 , n5577 );
and ( n11445 , n11443 , n11444 );
or ( n11446 , n11351 , n11445 );
xnor ( n11447 , n4073 , n5529 );
and ( n11448 , n11446 , n11447 );
or ( n11449 , n11349 , n11448 );
xnor ( n11450 , n4063 , n5526 );
and ( n11451 , n11449 , n11450 );
or ( n11452 , n11347 , n11451 );
xnor ( n11453 , n4053 , n5523 );
and ( n11454 , n11452 , n11453 );
or ( n11455 , n11345 , n11454 );
xnor ( n11456 , n4043 , n5520 );
and ( n11457 , n11455 , n11456 );
or ( n11458 , n11343 , n11457 );
xnor ( n11459 , n4033 , n5517 );
and ( n11460 , n11458 , n11459 );
or ( n11461 , n11341 , n11460 );
xnor ( n11462 , n4023 , n5514 );
and ( n11463 , n11461 , n11462 );
or ( n11464 , n11339 , n11463 );
xnor ( n11465 , n4013 , n5511 );
and ( n11466 , n11464 , n11465 );
or ( n11467 , n11337 , n11466 );
xnor ( n11468 , n4003 , n5508 );
and ( n11469 , n11467 , n11468 );
or ( n11470 , n11335 , n11469 );
xnor ( n11471 , n3993 , n5505 );
and ( n11472 , n11470 , n11471 );
or ( n11473 , n11333 , n11472 );
xnor ( n11474 , n3983 , n5502 );
and ( n11475 , n11473 , n11474 );
or ( n11476 , n11331 , n11475 );
xnor ( n11477 , n11327 , n5499 );
and ( n11478 , n11476 , n11477 );
or ( n11479 , n11329 , n11478 );
and ( n11480 , n11322 , n11479 );
not ( n11481 , n5496 );
and ( n11482 , n11481 , n11320 );
and ( n11483 , n11482 , n11321 );
or ( n11484 , n11480 , n11483 );
not ( n11485 , n11484 );
or ( n11486 , n11485 , n3290 );
and ( n11487 , n11486 , n3630 );
or ( n11488 , n11484 , n3290 );
and ( n11489 , n11488 , n3628 );
xor ( n11490 , n3770 , n5496 );
not ( n11491 , n11490 );
not ( n11492 , n5499 );
and ( n11493 , n11492 , n3819 );
not ( n11494 , n5502 );
and ( n11495 , n11494 , n3983 );
not ( n11496 , n5505 );
and ( n11497 , n11496 , n3993 );
not ( n11498 , n5508 );
and ( n11499 , n11498 , n4003 );
not ( n11500 , n5511 );
and ( n11501 , n11500 , n4013 );
not ( n11502 , n5514 );
and ( n11503 , n11502 , n4023 );
not ( n11504 , n5517 );
and ( n11505 , n11504 , n4033 );
not ( n11506 , n5520 );
and ( n11507 , n11506 , n4043 );
not ( n11508 , n5523 );
and ( n11509 , n11508 , n4053 );
not ( n11510 , n5526 );
and ( n11511 , n11510 , n4063 );
not ( n11512 , n5529 );
and ( n11513 , n11512 , n4073 );
not ( n11514 , n5577 );
and ( n11515 , n11514 , n4083 );
not ( n11516 , n5587 );
and ( n11517 , n11516 , n4093 );
not ( n11518 , n5597 );
and ( n11519 , n11518 , n4103 );
not ( n11520 , n5607 );
and ( n11521 , n11520 , n4113 );
not ( n11522 , n5617 );
and ( n11523 , n11522 , n4123 );
not ( n11524 , n5627 );
and ( n11525 , n11524 , n4133 );
not ( n11526 , n5637 );
and ( n11527 , n11526 , n4143 );
not ( n11528 , n5647 );
and ( n11529 , n11528 , n4153 );
not ( n11530 , n5657 );
and ( n11531 , n11530 , n4163 );
not ( n11532 , n5667 );
and ( n11533 , n11532 , n4173 );
not ( n11534 , n5677 );
and ( n11535 , n11534 , n4183 );
not ( n11536 , n5687 );
and ( n11537 , n11536 , n4193 );
not ( n11538 , n5697 );
and ( n11539 , n11538 , n4203 );
not ( n11540 , n5707 );
and ( n11541 , n11540 , n4213 );
not ( n11542 , n5717 );
and ( n11543 , n11542 , n4223 );
not ( n11544 , n5727 );
and ( n11545 , n11544 , n4233 );
not ( n11546 , n5737 );
and ( n11547 , n11546 , n4243 );
not ( n11548 , n5747 );
and ( n11549 , n11548 , n4257 );
not ( n11550 , n5757 );
and ( n11551 , n11550 , n3785 );
not ( n11552 , n5492 );
and ( n11553 , n11552 , n3795 );
xnor ( n11554 , n3785 , n5757 );
and ( n11555 , n11553 , n11554 );
or ( n11556 , n11551 , n11555 );
xnor ( n11557 , n4257 , n5747 );
and ( n11558 , n11556 , n11557 );
or ( n11559 , n11549 , n11558 );
xnor ( n11560 , n4243 , n5737 );
and ( n11561 , n11559 , n11560 );
or ( n11562 , n11547 , n11561 );
xnor ( n11563 , n4233 , n5727 );
and ( n11564 , n11562 , n11563 );
or ( n11565 , n11545 , n11564 );
xnor ( n11566 , n4223 , n5717 );
and ( n11567 , n11565 , n11566 );
or ( n11568 , n11543 , n11567 );
xnor ( n11569 , n4213 , n5707 );
and ( n11570 , n11568 , n11569 );
or ( n11571 , n11541 , n11570 );
xnor ( n11572 , n4203 , n5697 );
and ( n11573 , n11571 , n11572 );
or ( n11574 , n11539 , n11573 );
xnor ( n11575 , n4193 , n5687 );
and ( n11576 , n11574 , n11575 );
or ( n11577 , n11537 , n11576 );
xnor ( n11578 , n4183 , n5677 );
and ( n11579 , n11577 , n11578 );
or ( n11580 , n11535 , n11579 );
xnor ( n11581 , n4173 , n5667 );
and ( n11582 , n11580 , n11581 );
or ( n11583 , n11533 , n11582 );
xnor ( n11584 , n4163 , n5657 );
and ( n11585 , n11583 , n11584 );
or ( n11586 , n11531 , n11585 );
xnor ( n11587 , n4153 , n5647 );
and ( n11588 , n11586 , n11587 );
or ( n11589 , n11529 , n11588 );
xnor ( n11590 , n4143 , n5637 );
and ( n11591 , n11589 , n11590 );
or ( n11592 , n11527 , n11591 );
xnor ( n11593 , n4133 , n5627 );
and ( n11594 , n11592 , n11593 );
or ( n11595 , n11525 , n11594 );
xnor ( n11596 , n4123 , n5617 );
and ( n11597 , n11595 , n11596 );
or ( n11598 , n11523 , n11597 );
xnor ( n11599 , n4113 , n5607 );
and ( n11600 , n11598 , n11599 );
or ( n11601 , n11521 , n11600 );
xnor ( n11602 , n4103 , n5597 );
and ( n11603 , n11601 , n11602 );
or ( n11604 , n11519 , n11603 );
xnor ( n11605 , n4093 , n5587 );
and ( n11606 , n11604 , n11605 );
or ( n11607 , n11517 , n11606 );
xnor ( n11608 , n4083 , n5577 );
and ( n11609 , n11607 , n11608 );
or ( n11610 , n11515 , n11609 );
xnor ( n11611 , n4073 , n5529 );
and ( n11612 , n11610 , n11611 );
or ( n11613 , n11513 , n11612 );
xnor ( n11614 , n4063 , n5526 );
and ( n11615 , n11613 , n11614 );
or ( n11616 , n11511 , n11615 );
xnor ( n11617 , n4053 , n5523 );
and ( n11618 , n11616 , n11617 );
or ( n11619 , n11509 , n11618 );
xnor ( n11620 , n4043 , n5520 );
and ( n11621 , n11619 , n11620 );
or ( n11622 , n11507 , n11621 );
xnor ( n11623 , n4033 , n5517 );
and ( n11624 , n11622 , n11623 );
or ( n11625 , n11505 , n11624 );
xnor ( n11626 , n4023 , n5514 );
and ( n11627 , n11625 , n11626 );
or ( n11628 , n11503 , n11627 );
xnor ( n11629 , n4013 , n5511 );
and ( n11630 , n11628 , n11629 );
or ( n11631 , n11501 , n11630 );
xnor ( n11632 , n4003 , n5508 );
and ( n11633 , n11631 , n11632 );
or ( n11634 , n11499 , n11633 );
xnor ( n11635 , n3993 , n5505 );
and ( n11636 , n11634 , n11635 );
or ( n11637 , n11497 , n11636 );
xnor ( n11638 , n3983 , n5502 );
and ( n11639 , n11637 , n11638 );
or ( n11640 , n11495 , n11639 );
xnor ( n11641 , n3819 , n5499 );
and ( n11642 , n11640 , n11641 );
or ( n11643 , n11493 , n11642 );
and ( n11644 , n11491 , n11643 );
not ( n11645 , n3770 );
and ( n11646 , n11645 , n5496 );
and ( n11647 , n11646 , n11490 );
or ( n11648 , n11644 , n11647 );
or ( n11649 , n11648 , n3290 );
and ( n11650 , n11649 , n3626 );
not ( n11651 , n11648 );
or ( n11652 , n11651 , n3290 );
and ( n11653 , n11652 , n5285 );
xor ( n11654 , n3770 , n5496 );
xor ( n11655 , n3819 , n5499 );
or ( n11656 , n11654 , n11655 );
xor ( n11657 , n3983 , n5502 );
or ( n11658 , n11656 , n11657 );
xor ( n11659 , n3993 , n5505 );
or ( n11660 , n11658 , n11659 );
xor ( n11661 , n4003 , n5508 );
or ( n11662 , n11660 , n11661 );
xor ( n11663 , n4013 , n5511 );
or ( n11664 , n11662 , n11663 );
xor ( n11665 , n4023 , n5514 );
or ( n11666 , n11664 , n11665 );
xor ( n11667 , n4033 , n5517 );
or ( n11668 , n11666 , n11667 );
xor ( n11669 , n4043 , n5520 );
or ( n11670 , n11668 , n11669 );
xor ( n11671 , n4053 , n5523 );
or ( n11672 , n11670 , n11671 );
xor ( n11673 , n4063 , n5526 );
or ( n11674 , n11672 , n11673 );
xor ( n11675 , n4073 , n5529 );
or ( n11676 , n11674 , n11675 );
xor ( n11677 , n4083 , n5577 );
or ( n11678 , n11676 , n11677 );
xor ( n11679 , n4093 , n5587 );
or ( n11680 , n11678 , n11679 );
xor ( n11681 , n4103 , n5597 );
or ( n11682 , n11680 , n11681 );
xor ( n11683 , n4113 , n5607 );
or ( n11684 , n11682 , n11683 );
xor ( n11685 , n4123 , n5617 );
or ( n11686 , n11684 , n11685 );
xor ( n11687 , n4133 , n5627 );
or ( n11688 , n11686 , n11687 );
xor ( n11689 , n4143 , n5637 );
or ( n11690 , n11688 , n11689 );
xor ( n11691 , n4153 , n5647 );
or ( n11692 , n11690 , n11691 );
xor ( n11693 , n4163 , n5657 );
or ( n11694 , n11692 , n11693 );
xor ( n11695 , n4173 , n5667 );
or ( n11696 , n11694 , n11695 );
xor ( n11697 , n4183 , n5677 );
or ( n11698 , n11696 , n11697 );
xor ( n11699 , n4193 , n5687 );
or ( n11700 , n11698 , n11699 );
xor ( n11701 , n4203 , n5697 );
or ( n11702 , n11700 , n11701 );
xor ( n11703 , n4213 , n5707 );
or ( n11704 , n11702 , n11703 );
xor ( n11705 , n4223 , n5717 );
or ( n11706 , n11704 , n11705 );
xor ( n11707 , n4233 , n5727 );
or ( n11708 , n11706 , n11707 );
xor ( n11709 , n4243 , n5737 );
or ( n11710 , n11708 , n11709 );
xor ( n11711 , n4257 , n5747 );
or ( n11712 , n11710 , n11711 );
xor ( n11713 , n3785 , n5757 );
or ( n11714 , n11712 , n11713 );
xor ( n11715 , n3795 , n5492 );
or ( n11716 , n11714 , n11715 );
not ( n11717 , n11716 );
not ( n11718 , n11717 );
or ( n11719 , n11718 , n3290 );
and ( n11720 , n11719 , n6217 );
or ( n11721 , n11717 , n3290 );
and ( n11722 , n11721 , n6709 );
xor ( n11723 , n3770 , n5496 );
not ( n11724 , n11723 );
not ( n11725 , n3819 );
and ( n11726 , n11725 , n5499 );
not ( n11727 , n3983 );
and ( n11728 , n11727 , n5502 );
not ( n11729 , n3993 );
and ( n11730 , n11729 , n5505 );
not ( n11731 , n4003 );
and ( n11732 , n11731 , n5508 );
not ( n11733 , n4013 );
and ( n11734 , n11733 , n5511 );
not ( n11735 , n4023 );
and ( n11736 , n11735 , n5514 );
not ( n11737 , n4033 );
and ( n11738 , n11737 , n5517 );
not ( n11739 , n4043 );
and ( n11740 , n11739 , n5520 );
not ( n11741 , n4053 );
and ( n11742 , n11741 , n5523 );
not ( n11743 , n4063 );
and ( n11744 , n11743 , n5526 );
not ( n11745 , n4073 );
and ( n11746 , n11745 , n5529 );
not ( n11747 , n4083 );
and ( n11748 , n11747 , n5577 );
not ( n11749 , n4093 );
and ( n11750 , n11749 , n5587 );
not ( n11751 , n4103 );
and ( n11752 , n11751 , n5597 );
not ( n11753 , n4113 );
and ( n11754 , n11753 , n5607 );
not ( n11755 , n4123 );
and ( n11756 , n11755 , n5617 );
not ( n11757 , n4133 );
and ( n11758 , n11757 , n5627 );
not ( n11759 , n4143 );
and ( n11760 , n11759 , n5637 );
not ( n11761 , n4153 );
and ( n11762 , n11761 , n5647 );
not ( n11763 , n4163 );
and ( n11764 , n11763 , n5657 );
not ( n11765 , n4173 );
and ( n11766 , n11765 , n5667 );
not ( n11767 , n4183 );
and ( n11768 , n11767 , n5677 );
not ( n11769 , n4193 );
and ( n11770 , n11769 , n5687 );
not ( n11771 , n4203 );
and ( n11772 , n11771 , n5697 );
not ( n11773 , n4213 );
and ( n11774 , n11773 , n5707 );
not ( n11775 , n4223 );
and ( n11776 , n11775 , n5717 );
not ( n11777 , n4233 );
and ( n11778 , n11777 , n5727 );
not ( n11779 , n4243 );
and ( n11780 , n11779 , n5737 );
not ( n11781 , n4257 );
and ( n11782 , n11781 , n5747 );
not ( n11783 , n3785 );
and ( n11784 , n11783 , n5757 );
not ( n11785 , n3795 );
and ( n11786 , n11785 , n5492 );
xnor ( n11787 , n3785 , n5757 );
and ( n11788 , n11786 , n11787 );
or ( n11789 , n11784 , n11788 );
xnor ( n11790 , n4257 , n5747 );
and ( n11791 , n11789 , n11790 );
or ( n11792 , n11782 , n11791 );
xnor ( n11793 , n4243 , n5737 );
and ( n11794 , n11792 , n11793 );
or ( n11795 , n11780 , n11794 );
xnor ( n11796 , n4233 , n5727 );
and ( n11797 , n11795 , n11796 );
or ( n11798 , n11778 , n11797 );
xnor ( n11799 , n4223 , n5717 );
and ( n11800 , n11798 , n11799 );
or ( n11801 , n11776 , n11800 );
xnor ( n11802 , n4213 , n5707 );
and ( n11803 , n11801 , n11802 );
or ( n11804 , n11774 , n11803 );
xnor ( n11805 , n4203 , n5697 );
and ( n11806 , n11804 , n11805 );
or ( n11807 , n11772 , n11806 );
xnor ( n11808 , n4193 , n5687 );
and ( n11809 , n11807 , n11808 );
or ( n11810 , n11770 , n11809 );
xnor ( n11811 , n4183 , n5677 );
and ( n11812 , n11810 , n11811 );
or ( n11813 , n11768 , n11812 );
xnor ( n11814 , n4173 , n5667 );
and ( n11815 , n11813 , n11814 );
or ( n11816 , n11766 , n11815 );
xnor ( n11817 , n4163 , n5657 );
and ( n11818 , n11816 , n11817 );
or ( n11819 , n11764 , n11818 );
xnor ( n11820 , n4153 , n5647 );
and ( n11821 , n11819 , n11820 );
or ( n11822 , n11762 , n11821 );
xnor ( n11823 , n4143 , n5637 );
and ( n11824 , n11822 , n11823 );
or ( n11825 , n11760 , n11824 );
xnor ( n11826 , n4133 , n5627 );
and ( n11827 , n11825 , n11826 );
or ( n11828 , n11758 , n11827 );
xnor ( n11829 , n4123 , n5617 );
and ( n11830 , n11828 , n11829 );
or ( n11831 , n11756 , n11830 );
xnor ( n11832 , n4113 , n5607 );
and ( n11833 , n11831 , n11832 );
or ( n11834 , n11754 , n11833 );
xnor ( n11835 , n4103 , n5597 );
and ( n11836 , n11834 , n11835 );
or ( n11837 , n11752 , n11836 );
xnor ( n11838 , n4093 , n5587 );
and ( n11839 , n11837 , n11838 );
or ( n11840 , n11750 , n11839 );
xnor ( n11841 , n4083 , n5577 );
and ( n11842 , n11840 , n11841 );
or ( n11843 , n11748 , n11842 );
xnor ( n11844 , n4073 , n5529 );
and ( n11845 , n11843 , n11844 );
or ( n11846 , n11746 , n11845 );
xnor ( n11847 , n4063 , n5526 );
and ( n11848 , n11846 , n11847 );
or ( n11849 , n11744 , n11848 );
xnor ( n11850 , n4053 , n5523 );
and ( n11851 , n11849 , n11850 );
or ( n11852 , n11742 , n11851 );
xnor ( n11853 , n4043 , n5520 );
and ( n11854 , n11852 , n11853 );
or ( n11855 , n11740 , n11854 );
xnor ( n11856 , n4033 , n5517 );
and ( n11857 , n11855 , n11856 );
or ( n11858 , n11738 , n11857 );
xnor ( n11859 , n4023 , n5514 );
and ( n11860 , n11858 , n11859 );
or ( n11861 , n11736 , n11860 );
xnor ( n11862 , n4013 , n5511 );
and ( n11863 , n11861 , n11862 );
or ( n11864 , n11734 , n11863 );
xnor ( n11865 , n4003 , n5508 );
and ( n11866 , n11864 , n11865 );
or ( n11867 , n11732 , n11866 );
xnor ( n11868 , n3993 , n5505 );
and ( n11869 , n11867 , n11868 );
or ( n11870 , n11730 , n11869 );
xnor ( n11871 , n3983 , n5502 );
and ( n11872 , n11870 , n11871 );
or ( n11873 , n11728 , n11872 );
xnor ( n11874 , n3819 , n5499 );
and ( n11875 , n11873 , n11874 );
or ( n11876 , n11726 , n11875 );
and ( n11877 , n11724 , n11876 );
not ( n11878 , n5496 );
and ( n11879 , n11878 , n3770 );
and ( n11880 , n11879 , n11723 );
or ( n11881 , n11877 , n11880 );
not ( n11882 , n11881 );
or ( n11883 , n11882 , n3290 );
and ( n11884 , n11883 , n6215 );
or ( n11885 , n11881 , n3290 );
and ( n11886 , n11885 , n6707 );
and ( n11887 , n11485 , n6213 );
and ( n11888 , n11484 , n6212 );
and ( n11889 , n11648 , n6705 );
and ( n11890 , n11651 , n6704 );
and ( n11891 , n11718 , n6716 );
and ( n11892 , n11717 , n6715 );
and ( n11893 , n11882 , n6719 );
and ( n11894 , n11881 , n6724 );
or ( n11895 , n11487 , n11489 , n11650 , n11653 , n11720 , n11722 , n11884 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 );
and ( n11896 , n11895 , n3066 );
or ( n11897 , n11313 , n11896 );
and ( n11898 , n11897 , n2422 );
and ( n11899 , n3290 , n2428 );
or ( n11900 , n11898 , n11899 );
buf ( n11901 , n11900 );
buf ( n11902 , n2424 );
buf ( n11903 , n2281 );
buf ( n11904 , n2280 );
not ( n11905 , n3260 );
and ( n11906 , n3789 , n3631 );
and ( n11907 , n5156 , n5280 );
or ( n11908 , n5250 , n5188 );
buf ( n11909 , n11908 );
and ( n11910 , n3789 , n11909 );
or ( n11911 , n11907 , n11910 );
and ( n11912 , n11911 , n5285 );
and ( n11913 , n6207 , n5280 );
and ( n11914 , n3789 , n11909 );
or ( n11915 , n11913 , n11914 );
and ( n11916 , n11915 , n6218 );
and ( n11917 , n6700 , n5280 );
and ( n11918 , n3789 , n11909 );
or ( n11919 , n11917 , n11918 );
and ( n11920 , n11919 , n6710 );
and ( n11921 , n5492 , n5280 );
and ( n11922 , n3789 , n11909 );
or ( n11923 , n11921 , n11922 );
and ( n11924 , n11923 , n6717 );
and ( n11925 , n3363 , n6719 );
and ( n11926 , n5492 , n5280 );
and ( n11927 , n3789 , n11909 );
or ( n11928 , n11926 , n11927 );
and ( n11929 , n11928 , n6724 );
or ( n11930 , n11906 , n11912 , n11916 , n11920 , n11924 , n11925 , n11929 );
and ( n11931 , n11905 , n11930 );
and ( n11932 , n3789 , n3260 );
or ( n11933 , n11931 , n11932 );
and ( n11934 , n11933 , n2422 );
and ( n11935 , n3789 , n2428 );
or ( n11936 , n11934 , n11935 );
buf ( n11937 , n11936 );
buf ( n11938 , n2424 );
buf ( n11939 , n2281 );
buf ( n11940 , n2280 );
not ( n11941 , n3260 );
and ( n11942 , n3779 , n3631 );
and ( n11943 , n7043 , n5280 );
and ( n11944 , n3779 , n11909 );
or ( n11945 , n11943 , n11944 );
and ( n11946 , n11945 , n5285 );
and ( n11947 , n7054 , n5280 );
and ( n11948 , n3779 , n11909 );
or ( n11949 , n11947 , n11948 );
and ( n11950 , n11949 , n6218 );
and ( n11951 , n7065 , n5280 );
and ( n11952 , n3779 , n11909 );
or ( n11953 , n11951 , n11952 );
and ( n11954 , n11953 , n6710 );
and ( n11955 , n5757 , n5280 );
and ( n11956 , n3779 , n11909 );
or ( n11957 , n11955 , n11956 );
and ( n11958 , n11957 , n6717 );
and ( n11959 , n3776 , n6719 );
and ( n11960 , n7077 , n5280 );
and ( n11961 , n3779 , n11909 );
or ( n11962 , n11960 , n11961 );
and ( n11963 , n11962 , n6724 );
or ( n11964 , n11942 , n11946 , n11950 , n11954 , n11958 , n11959 , n11963 );
and ( n11965 , n11941 , n11964 );
and ( n11966 , n3779 , n3260 );
or ( n11967 , n11965 , n11966 );
and ( n11968 , n11967 , n2422 );
and ( n11969 , n3779 , n2428 );
or ( n11970 , n11968 , n11969 );
buf ( n11971 , n11970 );
buf ( n11972 , n2424 );
buf ( n11973 , n2281 );
buf ( n11974 , n2280 );
not ( n11975 , n3260 );
and ( n11976 , n4251 , n3631 );
and ( n11977 , n7117 , n5280 );
and ( n11978 , n4251 , n11909 );
or ( n11979 , n11977 , n11978 );
and ( n11980 , n11979 , n5285 );
and ( n11981 , n7128 , n5280 );
and ( n11982 , n4251 , n11909 );
or ( n11983 , n11981 , n11982 );
and ( n11984 , n11983 , n6218 );
and ( n11985 , n7139 , n5280 );
and ( n11986 , n4251 , n11909 );
or ( n11987 , n11985 , n11986 );
and ( n11988 , n11987 , n6710 );
and ( n11989 , n5747 , n5280 );
and ( n11990 , n4251 , n11909 );
or ( n11991 , n11989 , n11990 );
and ( n11992 , n11991 , n6717 );
and ( n11993 , n4249 , n6719 );
and ( n11994 , n7151 , n5280 );
and ( n11995 , n4251 , n11909 );
or ( n11996 , n11994 , n11995 );
and ( n11997 , n11996 , n6724 );
or ( n11998 , n11976 , n11980 , n11984 , n11988 , n11992 , n11993 , n11997 );
and ( n11999 , n11975 , n11998 );
and ( n12000 , n4251 , n3260 );
or ( n12001 , n11999 , n12000 );
and ( n12002 , n12001 , n2422 );
and ( n12003 , n4251 , n2428 );
or ( n12004 , n12002 , n12003 );
buf ( n12005 , n12004 );
buf ( n12006 , n2424 );
buf ( n12007 , n2281 );
buf ( n12008 , n2280 );
not ( n12009 , n3260 );
and ( n12010 , n4237 , n3631 );
and ( n12011 , n7191 , n5280 );
and ( n12012 , n4237 , n11909 );
or ( n12013 , n12011 , n12012 );
and ( n12014 , n12013 , n5285 );
and ( n12015 , n7202 , n5280 );
and ( n12016 , n4237 , n11909 );
or ( n12017 , n12015 , n12016 );
and ( n12018 , n12017 , n6218 );
and ( n12019 , n7213 , n5280 );
and ( n12020 , n4237 , n11909 );
or ( n12021 , n12019 , n12020 );
and ( n12022 , n12021 , n6710 );
and ( n12023 , n5737 , n5280 );
and ( n12024 , n4237 , n11909 );
or ( n12025 , n12023 , n12024 );
and ( n12026 , n12025 , n6717 );
and ( n12027 , n4235 , n6719 );
and ( n12028 , n7225 , n5280 );
and ( n12029 , n4237 , n11909 );
or ( n12030 , n12028 , n12029 );
and ( n12031 , n12030 , n6724 );
or ( n12032 , n12010 , n12014 , n12018 , n12022 , n12026 , n12027 , n12031 );
and ( n12033 , n12009 , n12032 );
and ( n12034 , n4237 , n3260 );
or ( n12035 , n12033 , n12034 );
and ( n12036 , n12035 , n2422 );
and ( n12037 , n4237 , n2428 );
or ( n12038 , n12036 , n12037 );
buf ( n12039 , n12038 );
buf ( n12040 , n2424 );
buf ( n12041 , n2281 );
buf ( n12042 , n2280 );
not ( n12043 , n3260 );
and ( n12044 , n4227 , n3631 );
and ( n12045 , n7265 , n5280 );
and ( n12046 , n4227 , n11909 );
or ( n12047 , n12045 , n12046 );
and ( n12048 , n12047 , n5285 );
and ( n12049 , n7276 , n5280 );
and ( n12050 , n4227 , n11909 );
or ( n12051 , n12049 , n12050 );
and ( n12052 , n12051 , n6218 );
and ( n12053 , n7287 , n5280 );
and ( n12054 , n4227 , n11909 );
or ( n12055 , n12053 , n12054 );
and ( n12056 , n12055 , n6710 );
and ( n12057 , n5727 , n5280 );
and ( n12058 , n4227 , n11909 );
or ( n12059 , n12057 , n12058 );
and ( n12060 , n12059 , n6717 );
and ( n12061 , n4225 , n6719 );
nand ( n12062 , n7299 , n5280 );
and ( n12063 , n4227 , n11909 );
or ( n12064 , n12062 , n12063 );
and ( n12065 , n12064 , n6724 );
or ( n12066 , n12044 , n12048 , n12052 , n12056 , n12060 , n12061 , n12065 );
and ( n12067 , n12043 , n12066 );
and ( n12068 , n4227 , n3260 );
or ( n12069 , n12067 , n12068 );
and ( n12070 , n12069 , n2422 );
and ( n12071 , n4227 , n2428 );
or ( n12072 , n12070 , n12071 );
buf ( n12073 , n12072 );
buf ( n12074 , n2424 );
buf ( n12075 , n2281 );
buf ( n12076 , n2280 );
not ( n12077 , n3260 );
and ( n12078 , n4217 , n3631 );
and ( n12079 , n7339 , n5280 );
and ( n12080 , n4217 , n11909 );
or ( n12081 , n12079 , n12080 );
and ( n12082 , n12081 , n5285 );
and ( n12083 , n7350 , n5280 );
and ( n12084 , n4217 , n11909 );
or ( n12085 , n12083 , n12084 );
and ( n12086 , n12085 , n6218 );
and ( n12087 , n7361 , n5280 );
and ( n12088 , n4217 , n11909 );
or ( n12089 , n12087 , n12088 );
and ( n12090 , n12089 , n6710 );
and ( n12091 , n5717 , n5280 );
and ( n12092 , n4217 , n11909 );
or ( n12093 , n12091 , n12092 );
and ( n12094 , n12093 , n6717 );
and ( n12095 , n4215 , n6719 );
and ( n12096 , n7373 , n5280 );
and ( n12097 , n4217 , n11909 );
or ( n12098 , n12096 , n12097 );
and ( n12099 , n12098 , n6724 );
or ( n12100 , n12078 , n12082 , n12086 , n12090 , n12094 , n12095 , n12099 );
and ( n12101 , n12077 , n12100 );
and ( n12102 , n4217 , n3260 );
or ( n12103 , n12101 , n12102 );
and ( n12104 , n12103 , n2422 );
and ( n12105 , n4217 , n2428 );
or ( n12106 , n12104 , n12105 );
buf ( n12107 , n12106 );
buf ( n12108 , n2424 );
buf ( n12109 , n2281 );
buf ( n12110 , n2280 );
not ( n12111 , n3260 );
and ( n12112 , n4207 , n3631 );
and ( n12113 , n7413 , n5280 );
and ( n12114 , n4207 , n11909 );
or ( n12115 , n12113 , n12114 );
and ( n12116 , n12115 , n5285 );
and ( n12117 , n7424 , n5280 );
and ( n12118 , n4207 , n11909 );
or ( n12119 , n12117 , n12118 );
and ( n12120 , n12119 , n6218 );
and ( n12121 , n7435 , n5280 );
and ( n12122 , n4207 , n11909 );
or ( n12123 , n12121 , n12122 );
and ( n12124 , n12123 , n6710 );
and ( n12125 , n5707 , n5280 );
and ( n12126 , n4207 , n11909 );
or ( n12127 , n12125 , n12126 );
and ( n12128 , n12127 , n6717 );
and ( n12129 , n4205 , n6719 );
and ( n12130 , n7447 , n5280 );
and ( n12131 , n4207 , n11909 );
or ( n12132 , n12130 , n12131 );
and ( n12133 , n12132 , n6724 );
or ( n12134 , n12112 , n12116 , n12120 , n12124 , n12128 , n12129 , n12133 );
and ( n12135 , n12111 , n12134 );
and ( n12136 , n4207 , n3260 );
or ( n12137 , n12135 , n12136 );
and ( n12138 , n12137 , n2422 );
and ( n12139 , n4207 , n2428 );
or ( n12140 , n12138 , n12139 );
buf ( n12141 , n12140 );
buf ( n12142 , n2424 );
buf ( n12143 , n2281 );
buf ( n12144 , n2280 );
not ( n12145 , n3260 );
and ( n12146 , n4197 , n3631 );
and ( n12147 , n7487 , n5280 );
and ( n12148 , n4197 , n11909 );
or ( n12149 , n12147 , n12148 );
and ( n12150 , n12149 , n5285 );
and ( n12151 , n7498 , n5280 );
and ( n12152 , n4197 , n11909 );
or ( n12153 , n12151 , n12152 );
and ( n12154 , n12153 , n6218 );
and ( n12155 , n7509 , n5280 );
and ( n12156 , n4197 , n11909 );
or ( n12157 , n12155 , n12156 );
and ( n12158 , n12157 , n6710 );
and ( n12159 , n5697 , n5280 );
and ( n12160 , n4197 , n11909 );
or ( n12161 , n12159 , n12160 );
and ( n12162 , n12161 , n6717 );
and ( n12163 , n4195 , n6719 );
and ( n12164 , n7521 , n5280 );
and ( n12165 , n4197 , n11909 );
or ( n12166 , n12164 , n12165 );
and ( n12167 , n12166 , n6724 );
or ( n12168 , n12146 , n12150 , n12154 , n12158 , n12162 , n12163 , n12167 );
and ( n12169 , n12145 , n12168 );
and ( n12170 , n4197 , n3260 );
or ( n12171 , n12169 , n12170 );
and ( n12172 , n12171 , n2422 );
and ( n12173 , n4197 , n2428 );
or ( n12174 , n12172 , n12173 );
buf ( n12175 , n12174 );
buf ( n12176 , n2424 );
buf ( n12177 , n2281 );
buf ( n12178 , n2280 );
not ( n12179 , n3260 );
and ( n12180 , n4187 , n3631 );
and ( n12181 , n7561 , n5280 );
and ( n12182 , n4187 , n11909 );
or ( n12183 , n12181 , n12182 );
and ( n12184 , n12183 , n5285 );
and ( n12185 , n7572 , n5280 );
and ( n12186 , n4187 , n11909 );
or ( n12187 , n12185 , n12186 );
and ( n12188 , n12187 , n6218 );
and ( n12189 , n7583 , n5280 );
and ( n12190 , n4187 , n11909 );
or ( n12191 , n12189 , n12190 );
and ( n12192 , n12191 , n6710 );
and ( n12193 , n5687 , n5280 );
and ( n12194 , n4187 , n11909 );
or ( n12195 , n12193 , n12194 );
and ( n12196 , n12195 , n6717 );
and ( n12197 , n4185 , n6719 );
and ( n12198 , n7595 , n5280 );
and ( n12199 , n4187 , n11909 );
or ( n12200 , n12198 , n12199 );
and ( n12201 , n12200 , n6724 );
or ( n12202 , n12180 , n12184 , n12188 , n12192 , n12196 , n12197 , n12201 );
and ( n12203 , n12179 , n12202 );
and ( n12204 , n4187 , n3260 );
or ( n12205 , n12203 , n12204 );
and ( n12206 , n12205 , n2422 );
and ( n12207 , n4187 , n2428 );
or ( n12208 , n12206 , n12207 );
buf ( n12209 , n12208 );
buf ( n12210 , n2424 );
buf ( n12211 , n2281 );
buf ( n12212 , n2280 );
not ( n12213 , n3260 );
and ( n12214 , n4177 , n3631 );
and ( n12215 , n7635 , n5280 );
and ( n12216 , n4177 , n11909 );
or ( n12217 , n12215 , n12216 );
and ( n12218 , n12217 , n5285 );
and ( n12219 , n7646 , n5280 );
and ( n12220 , n4177 , n11909 );
or ( n12221 , n12219 , n12220 );
and ( n12222 , n12221 , n6218 );
and ( n12223 , n7657 , n5280 );
and ( n12224 , n4177 , n11909 );
or ( n12225 , n12223 , n12224 );
and ( n12226 , n12225 , n6710 );
and ( n12227 , n5677 , n5280 );
and ( n12228 , n4177 , n11909 );
or ( n12229 , n12227 , n12228 );
and ( n12230 , n12229 , n6717 );
and ( n12231 , n4175 , n6719 );
and ( n12232 , n7669 , n5280 );
and ( n12233 , n4177 , n11909 );
or ( n12234 , n12232 , n12233 );
and ( n12235 , n12234 , n6724 );
or ( n12236 , n12214 , n12218 , n12222 , n12226 , n12230 , n12231 , n12235 );
and ( n12237 , n12213 , n12236 );
and ( n12238 , n4177 , n3260 );
or ( n12239 , n12237 , n12238 );
and ( n12240 , n12239 , n2422 );
and ( n12241 , n4177 , n2428 );
or ( n12242 , n12240 , n12241 );
buf ( n12243 , n12242 );
buf ( n12244 , n2424 );
buf ( n12245 , n2281 );
buf ( n12246 , n2280 );
not ( n12247 , n3260 );
and ( n12248 , n4167 , n3631 );
and ( n12249 , n7709 , n5280 );
and ( n12250 , n4167 , n11909 );
or ( n12251 , n12249 , n12250 );
and ( n12252 , n12251 , n5285 );
and ( n12253 , n7720 , n5280 );
and ( n12254 , n4167 , n11909 );
or ( n12255 , n12253 , n12254 );
and ( n12256 , n12255 , n6218 );
and ( n12257 , n7731 , n5280 );
and ( n12258 , n4167 , n11909 );
or ( n12259 , n12257 , n12258 );
and ( n12260 , n12259 , n6710 );
and ( n12261 , n5667 , n5280 );
and ( n12262 , n4167 , n11909 );
or ( n12263 , n12261 , n12262 );
and ( n12264 , n12263 , n6717 );
and ( n12265 , n4165 , n6719 );
and ( n12266 , n7743 , n5280 );
and ( n12267 , n4167 , n11909 );
or ( n12268 , n12266 , n12267 );
and ( n12269 , n12268 , n6724 );
or ( n12270 , n12248 , n12252 , n12256 , n12260 , n12264 , n12265 , n12269 );
and ( n12271 , n12247 , n12270 );
and ( n12272 , n4167 , n3260 );
or ( n12273 , n12271 , n12272 );
and ( n12274 , n12273 , n2422 );
and ( n12275 , n4167 , n2428 );
or ( n12276 , n12274 , n12275 );
buf ( n12277 , n12276 );
buf ( n12278 , n2424 );
buf ( n12279 , n2281 );
buf ( n12280 , n2280 );
not ( n12281 , n3260 );
and ( n12282 , n4157 , n3631 );
and ( n12283 , n7783 , n5280 );
and ( n12284 , n4157 , n11909 );
or ( n12285 , n12283 , n12284 );
and ( n12286 , n12285 , n5285 );
and ( n12287 , n7794 , n5280 );
and ( n12288 , n4157 , n11909 );
or ( n12289 , n12287 , n12288 );
and ( n12290 , n12289 , n6218 );
and ( n12291 , n7805 , n5280 );
and ( n12292 , n4157 , n11909 );
or ( n12293 , n12291 , n12292 );
and ( n12294 , n12293 , n6710 );
and ( n12295 , n5657 , n5280 );
and ( n12296 , n4157 , n11909 );
or ( n12297 , n12295 , n12296 );
and ( n12298 , n12297 , n6717 );
and ( n12299 , n4155 , n6719 );
and ( n12300 , n7817 , n5280 );
and ( n12301 , n4157 , n11909 );
or ( n12302 , n12300 , n12301 );
and ( n12303 , n12302 , n6724 );
or ( n12304 , n12282 , n12286 , n12290 , n12294 , n12298 , n12299 , n12303 );
and ( n12305 , n12281 , n12304 );
and ( n12306 , n4157 , n3260 );
or ( n12307 , n12305 , n12306 );
and ( n12308 , n12307 , n2422 );
and ( n12309 , n4157 , n2428 );
or ( n12310 , n12308 , n12309 );
buf ( n12311 , n12310 );
buf ( n12312 , n2424 );
buf ( n12313 , n2281 );
buf ( n12314 , n2280 );
not ( n12315 , n3260 );
and ( n12316 , n4147 , n3631 );
and ( n12317 , n7857 , n5280 );
and ( n12318 , n4147 , n11909 );
or ( n12319 , n12317 , n12318 );
and ( n12320 , n12319 , n5285 );
and ( n12321 , n7868 , n5280 );
and ( n12322 , n4147 , n11909 );
or ( n12323 , n12321 , n12322 );
and ( n12324 , n12323 , n6218 );
and ( n12325 , n7879 , n5280 );
and ( n12326 , n4147 , n11909 );
or ( n12327 , n12325 , n12326 );
and ( n12328 , n12327 , n6710 );
and ( n12329 , n5647 , n5280 );
and ( n12330 , n4147 , n11909 );
or ( n12331 , n12329 , n12330 );
and ( n12332 , n12331 , n6717 );
and ( n12333 , n4145 , n6719 );
and ( n12334 , n7891 , n5280 );
and ( n12335 , n4147 , n11909 );
or ( n12336 , n12334 , n12335 );
and ( n12337 , n12336 , n6724 );
or ( n12338 , n12316 , n12320 , n12324 , n12328 , n12332 , n12333 , n12337 );
and ( n12339 , n12315 , n12338 );
and ( n12340 , n4147 , n3260 );
or ( n12341 , n12339 , n12340 );
and ( n12342 , n12341 , n2422 );
and ( n12343 , n4147 , n2428 );
or ( n12344 , n12342 , n12343 );
buf ( n12345 , n12344 );
buf ( n12346 , n2424 );
buf ( n12347 , n2281 );
buf ( n12348 , n2280 );
not ( n12349 , n3260 );
and ( n12350 , n4137 , n3631 );
and ( n12351 , n7931 , n5280 );
and ( n12352 , n4137 , n11909 );
or ( n12353 , n12351 , n12352 );
and ( n12354 , n12353 , n5285 );
and ( n12355 , n7942 , n5280 );
and ( n12356 , n4137 , n11909 );
or ( n12357 , n12355 , n12356 );
and ( n12358 , n12357 , n6218 );
and ( n12359 , n7953 , n5280 );
and ( n12360 , n4137 , n11909 );
or ( n12361 , n12359 , n12360 );
and ( n12362 , n12361 , n6710 );
and ( n12363 , n5637 , n5280 );
and ( n12364 , n4137 , n11909 );
or ( n12365 , n12363 , n12364 );
and ( n12366 , n12365 , n6717 );
and ( n12367 , n4135 , n6719 );
and ( n12368 , n7965 , n5280 );
and ( n12369 , n4137 , n11909 );
or ( n12370 , n12368 , n12369 );
and ( n12371 , n12370 , n6724 );
or ( n12372 , n12350 , n12354 , n12358 , n12362 , n12366 , n12367 , n12371 );
and ( n12373 , n12349 , n12372 );
and ( n12374 , n4137 , n3260 );
or ( n12375 , n12373 , n12374 );
and ( n12376 , n12375 , n2422 );
and ( n12377 , n4137 , n2428 );
or ( n12378 , n12376 , n12377 );
buf ( n12379 , n12378 );
buf ( n12380 , n2424 );
buf ( n12381 , n2281 );
buf ( n12382 , n2280 );
not ( n12383 , n3260 );
and ( n12384 , n4127 , n3631 );
and ( n12385 , n8005 , n5280 );
and ( n12386 , n4127 , n11909 );
or ( n12387 , n12385 , n12386 );
and ( n12388 , n12387 , n5285 );
and ( n12389 , n8016 , n5280 );
and ( n12390 , n4127 , n11909 );
or ( n12391 , n12389 , n12390 );
and ( n12392 , n12391 , n6218 );
and ( n12393 , n8027 , n5280 );
and ( n12394 , n4127 , n11909 );
or ( n12395 , n12393 , n12394 );
and ( n12396 , n12395 , n6710 );
and ( n12397 , n5627 , n5280 );
and ( n12398 , n4127 , n11909 );
or ( n12399 , n12397 , n12398 );
and ( n12400 , n12399 , n6717 );
and ( n12401 , n4125 , n6719 );
and ( n12402 , n8039 , n5280 );
and ( n12403 , n4127 , n11909 );
or ( n12404 , n12402 , n12403 );
and ( n12405 , n12404 , n6724 );
or ( n12406 , n12384 , n12388 , n12392 , n12396 , n12400 , n12401 , n12405 );
and ( n12407 , n12383 , n12406 );
and ( n12408 , n4127 , n3260 );
or ( n12409 , n12407 , n12408 );
and ( n12410 , n12409 , n2422 );
and ( n12411 , n4127 , n2428 );
or ( n12412 , n12410 , n12411 );
buf ( n12413 , n12412 );
buf ( n12414 , n2424 );
buf ( n12415 , n2281 );
buf ( n12416 , n2280 );
not ( n12417 , n3260 );
and ( n12418 , n4117 , n3631 );
and ( n12419 , n8079 , n5280 );
and ( n12420 , n4117 , n11909 );
or ( n12421 , n12419 , n12420 );
and ( n12422 , n12421 , n5285 );
and ( n12423 , n8090 , n5280 );
and ( n12424 , n4117 , n11909 );
or ( n12425 , n12423 , n12424 );
and ( n12426 , n12425 , n6218 );
and ( n12427 , n8101 , n5280 );
and ( n12428 , n4117 , n11909 );
or ( n12429 , n12427 , n12428 );
and ( n12430 , n12429 , n6710 );
and ( n12431 , n5617 , n5280 );
and ( n12432 , n4117 , n11909 );
or ( n12433 , n12431 , n12432 );
and ( n12434 , n12433 , n6717 );
and ( n12435 , n4115 , n6719 );
and ( n12436 , n8113 , n5280 );
and ( n12437 , n4117 , n11909 );
or ( n12438 , n12436 , n12437 );
and ( n12439 , n12438 , n6724 );
or ( n12440 , n12418 , n12422 , n12426 , n12430 , n12434 , n12435 , n12439 );
and ( n12441 , n12417 , n12440 );
and ( n12442 , n4117 , n3260 );
or ( n12443 , n12441 , n12442 );
and ( n12444 , n12443 , n2422 );
and ( n12445 , n4117 , n2428 );
or ( n12446 , n12444 , n12445 );
buf ( n12447 , n12446 );
buf ( n12448 , n2424 );
buf ( n12449 , n2281 );
buf ( n12450 , n2280 );
not ( n12451 , n3260 );
and ( n12452 , n4107 , n3631 );
and ( n12453 , n8153 , n5280 );
and ( n12454 , n4107 , n11909 );
or ( n12455 , n12453 , n12454 );
and ( n12456 , n12455 , n5285 );
and ( n12457 , n8164 , n5280 );
and ( n12458 , n4107 , n11909 );
or ( n12459 , n12457 , n12458 );
and ( n12460 , n12459 , n6218 );
and ( n12461 , n8175 , n5280 );
and ( n12462 , n4107 , n11909 );
or ( n12463 , n12461 , n12462 );
and ( n12464 , n12463 , n6710 );
and ( n12465 , n5607 , n5280 );
and ( n12466 , n4107 , n11909 );
or ( n12467 , n12465 , n12466 );
and ( n12468 , n12467 , n6717 );
and ( n12469 , n4105 , n6719 );
and ( n12470 , n8187 , n5280 );
and ( n12471 , n4107 , n11909 );
or ( n12472 , n12470 , n12471 );
and ( n12473 , n12472 , n6724 );
or ( n12474 , n12452 , n12456 , n12460 , n12464 , n12468 , n12469 , n12473 );
and ( n12475 , n12451 , n12474 );
and ( n12476 , n4107 , n3260 );
or ( n12477 , n12475 , n12476 );
and ( n12478 , n12477 , n2422 );
and ( n12479 , n4107 , n2428 );
or ( n12480 , n12478 , n12479 );
buf ( n12481 , n12480 );
buf ( n12482 , n2424 );
buf ( n12483 , n2281 );
buf ( n12484 , n2280 );
not ( n12485 , n3260 );
and ( n12486 , n4097 , n3631 );
and ( n12487 , n8227 , n5280 );
and ( n12488 , n4097 , n11909 );
or ( n12489 , n12487 , n12488 );
and ( n12490 , n12489 , n5285 );
and ( n12491 , n8238 , n5280 );
and ( n12492 , n4097 , n11909 );
or ( n12493 , n12491 , n12492 );
and ( n12494 , n12493 , n6218 );
and ( n12495 , n8249 , n5280 );
and ( n12496 , n4097 , n11909 );
or ( n12497 , n12495 , n12496 );
and ( n12498 , n12497 , n6710 );
and ( n12499 , n5597 , n5280 );
and ( n12500 , n4097 , n11909 );
or ( n12501 , n12499 , n12500 );
and ( n12502 , n12501 , n6717 );
and ( n12503 , n4095 , n6719 );
and ( n12504 , n8261 , n5280 );
and ( n12505 , n4097 , n11909 );
or ( n12506 , n12504 , n12505 );
and ( n12507 , n12506 , n6724 );
or ( n12508 , n12486 , n12490 , n12494 , n12498 , n12502 , n12503 , n12507 );
and ( n12509 , n12485 , n12508 );
and ( n12510 , n4097 , n3260 );
or ( n12511 , n12509 , n12510 );
and ( n12512 , n12511 , n2422 );
and ( n12513 , n4097 , n2428 );
or ( n12514 , n12512 , n12513 );
buf ( n12515 , n12514 );
buf ( n12516 , n2424 );
buf ( n12517 , n2281 );
buf ( n12518 , n2280 );
not ( n12519 , n3260 );
and ( n12520 , n4087 , n3631 );
and ( n12521 , n8301 , n5280 );
and ( n12522 , n4087 , n11909 );
or ( n12523 , n12521 , n12522 );
and ( n12524 , n12523 , n5285 );
and ( n12525 , n8312 , n5280 );
and ( n12526 , n4087 , n11909 );
or ( n12527 , n12525 , n12526 );
and ( n12528 , n12527 , n6218 );
and ( n12529 , n8323 , n5280 );
and ( n12530 , n4087 , n11909 );
or ( n12531 , n12529 , n12530 );
and ( n12532 , n12531 , n6710 );
and ( n12533 , n5587 , n5280 );
and ( n12534 , n4087 , n11909 );
or ( n12535 , n12533 , n12534 );
and ( n12536 , n12535 , n6717 );
and ( n12537 , n4085 , n6719 );
and ( n12538 , n8335 , n5280 );
and ( n12539 , n4087 , n11909 );
or ( n12540 , n12538 , n12539 );
and ( n12541 , n12540 , n6724 );
or ( n12542 , n12520 , n12524 , n12528 , n12532 , n12536 , n12537 , n12541 );
and ( n12543 , n12519 , n12542 );
and ( n12544 , n4087 , n3260 );
or ( n12545 , n12543 , n12544 );
and ( n12546 , n12545 , n2422 );
and ( n12547 , n4087 , n2428 );
or ( n12548 , n12546 , n12547 );
buf ( n12549 , n12548 );
buf ( n12550 , n2424 );
buf ( n12551 , n2281 );
buf ( n12552 , n2280 );
not ( n12553 , n3260 );
and ( n12554 , n4077 , n3631 );
and ( n12555 , n8375 , n5280 );
and ( n12556 , n4077 , n11909 );
or ( n12557 , n12555 , n12556 );
and ( n12558 , n12557 , n5285 );
and ( n12559 , n8386 , n5280 );
and ( n12560 , n4077 , n11909 );
or ( n12561 , n12559 , n12560 );
and ( n12562 , n12561 , n6218 );
and ( n12563 , n8397 , n5280 );
and ( n12564 , n4077 , n11909 );
or ( n12565 , n12563 , n12564 );
and ( n12566 , n12565 , n6710 );
and ( n12567 , n5577 , n5280 );
and ( n12568 , n4077 , n11909 );
or ( n12569 , n12567 , n12568 );
and ( n12570 , n12569 , n6717 );
and ( n12571 , n4075 , n6719 );
and ( n12572 , n8409 , n5280 );
and ( n12573 , n4077 , n11909 );
or ( n12574 , n12572 , n12573 );
and ( n12575 , n12574 , n6724 );
or ( n12576 , n12554 , n12558 , n12562 , n12566 , n12570 , n12571 , n12575 );
and ( n12577 , n12553 , n12576 );
and ( n12578 , n4077 , n3260 );
or ( n12579 , n12577 , n12578 );
and ( n12580 , n12579 , n2422 );
and ( n12581 , n4077 , n2428 );
or ( n12582 , n12580 , n12581 );
buf ( n12583 , n12582 );
buf ( n12584 , n2424 );
buf ( n12585 , n2281 );
buf ( n12586 , n2280 );
not ( n12587 , n3260 );
and ( n12588 , n4067 , n3631 );
and ( n12589 , n8449 , n5280 );
and ( n12590 , n4067 , n11909 );
or ( n12591 , n12589 , n12590 );
and ( n12592 , n12591 , n5285 );
and ( n12593 , n8460 , n5280 );
and ( n12594 , n4067 , n11909 );
or ( n12595 , n12593 , n12594 );
and ( n12596 , n12595 , n6218 );
and ( n12597 , n8471 , n5280 );
and ( n12598 , n4067 , n11909 );
or ( n12599 , n12597 , n12598 );
and ( n12600 , n12599 , n6710 );
and ( n12601 , n5529 , n5280 );
and ( n12602 , n4067 , n11909 );
or ( n12603 , n12601 , n12602 );
and ( n12604 , n12603 , n6717 );
and ( n12605 , n4065 , n6719 );
and ( n12606 , n8483 , n5280 );
and ( n12607 , n4067 , n11909 );
or ( n12608 , n12606 , n12607 );
and ( n12609 , n12608 , n6724 );
or ( n12610 , n12588 , n12592 , n12596 , n12600 , n12604 , n12605 , n12609 );
and ( n12611 , n12587 , n12610 );
and ( n12612 , n4067 , n3260 );
or ( n12613 , n12611 , n12612 );
and ( n12614 , n12613 , n2422 );
and ( n12615 , n4067 , n2428 );
or ( n12616 , n12614 , n12615 );
buf ( n12617 , n12616 );
buf ( n12618 , n2424 );
buf ( n12619 , n2281 );
buf ( n12620 , n2280 );
not ( n12621 , n3260 );
and ( n12622 , n4057 , n3631 );
and ( n12623 , n8523 , n5280 );
and ( n12624 , n4057 , n11909 );
or ( n12625 , n12623 , n12624 );
and ( n12626 , n12625 , n5285 );
and ( n12627 , n8534 , n5280 );
and ( n12628 , n4057 , n11909 );
or ( n12629 , n12627 , n12628 );
and ( n12630 , n12629 , n6218 );
and ( n12631 , n8545 , n5280 );
and ( n12632 , n4057 , n11909 );
or ( n12633 , n12631 , n12632 );
and ( n12634 , n12633 , n6710 );
and ( n12635 , n5526 , n5280 );
and ( n12636 , n4057 , n11909 );
or ( n12637 , n12635 , n12636 );
and ( n12638 , n12637 , n6717 );
and ( n12639 , n4055 , n6719 );
and ( n12640 , n8557 , n5280 );
and ( n12641 , n4057 , n11909 );
or ( n12642 , n12640 , n12641 );
and ( n12643 , n12642 , n6724 );
or ( n12644 , n12622 , n12626 , n12630 , n12634 , n12638 , n12639 , n12643 );
and ( n12645 , n12621 , n12644 );
and ( n12646 , n4057 , n3260 );
or ( n12647 , n12645 , n12646 );
and ( n12648 , n12647 , n2422 );
and ( n12649 , n4057 , n2428 );
or ( n12650 , n12648 , n12649 );
buf ( n12651 , n12650 );
buf ( n12652 , n2424 );
buf ( n12653 , n2281 );
buf ( n12654 , n2280 );
not ( n12655 , n3260 );
and ( n12656 , n4047 , n3631 );
and ( n12657 , n8597 , n5280 );
and ( n12658 , n4047 , n11909 );
or ( n12659 , n12657 , n12658 );
and ( n12660 , n12659 , n5285 );
and ( n12661 , n8608 , n5280 );
and ( n12662 , n4047 , n11909 );
or ( n12663 , n12661 , n12662 );
and ( n12664 , n12663 , n6218 );
and ( n12665 , n8619 , n5280 );
and ( n12666 , n4047 , n11909 );
or ( n12667 , n12665 , n12666 );
and ( n12668 , n12667 , n6710 );
and ( n12669 , n5523 , n5280 );
and ( n12670 , n4047 , n11909 );
or ( n12671 , n12669 , n12670 );
and ( n12672 , n12671 , n6717 );
and ( n12673 , n4045 , n6719 );
and ( n12674 , n8631 , n5280 );
and ( n12675 , n4047 , n11909 );
or ( n12676 , n12674 , n12675 );
and ( n12677 , n12676 , n6724 );
or ( n12678 , n12656 , n12660 , n12664 , n12668 , n12672 , n12673 , n12677 );
and ( n12679 , n12655 , n12678 );
and ( n12680 , n4047 , n3260 );
or ( n12681 , n12679 , n12680 );
and ( n12682 , n12681 , n2422 );
and ( n12683 , n4047 , n2428 );
or ( n12684 , n12682 , n12683 );
buf ( n12685 , n12684 );
buf ( n12686 , n2424 );
buf ( n12687 , n2281 );
buf ( n12688 , n2280 );
not ( n12689 , n3260 );
and ( n12690 , n4037 , n3631 );
and ( n12691 , n8671 , n5280 );
and ( n12692 , n4037 , n11909 );
or ( n12693 , n12691 , n12692 );
and ( n12694 , n12693 , n5285 );
and ( n12695 , n8682 , n5280 );
and ( n12696 , n4037 , n11909 );
or ( n12697 , n12695 , n12696 );
and ( n12698 , n12697 , n6218 );
and ( n12699 , n8693 , n5280 );
and ( n12700 , n4037 , n11909 );
or ( n12701 , n12699 , n12700 );
and ( n12702 , n12701 , n6710 );
and ( n12703 , n5520 , n5280 );
and ( n12704 , n4037 , n11909 );
or ( n12705 , n12703 , n12704 );
and ( n12706 , n12705 , n6717 );
and ( n12707 , n4035 , n6719 );
and ( n12708 , n8705 , n5280 );
and ( n12709 , n4037 , n11909 );
or ( n12710 , n12708 , n12709 );
and ( n12711 , n12710 , n6724 );
or ( n12712 , n12690 , n12694 , n12698 , n12702 , n12706 , n12707 , n12711 );
and ( n12713 , n12689 , n12712 );
and ( n12714 , n4037 , n3260 );
or ( n12715 , n12713 , n12714 );
and ( n12716 , n12715 , n2422 );
and ( n12717 , n4037 , n2428 );
or ( n12718 , n12716 , n12717 );
buf ( n12719 , n12718 );
buf ( n12720 , n2424 );
buf ( n12721 , n2281 );
buf ( n12722 , n2280 );
not ( n12723 , n3260 );
and ( n12724 , n4027 , n3631 );
and ( n12725 , n8745 , n5280 );
and ( n12726 , n4027 , n11909 );
or ( n12727 , n12725 , n12726 );
and ( n12728 , n12727 , n5285 );
and ( n12729 , n8756 , n5280 );
and ( n12730 , n4027 , n11909 );
or ( n12731 , n12729 , n12730 );
and ( n12732 , n12731 , n6218 );
and ( n12733 , n8767 , n5280 );
and ( n12734 , n4027 , n11909 );
or ( n12735 , n12733 , n12734 );
and ( n12736 , n12735 , n6710 );
and ( n12737 , n5517 , n5280 );
and ( n12738 , n4027 , n11909 );
or ( n12739 , n12737 , n12738 );
and ( n12740 , n12739 , n6717 );
and ( n12741 , n4025 , n6719 );
and ( n12742 , n8779 , n5280 );
and ( n12743 , n4027 , n11909 );
or ( n12744 , n12742 , n12743 );
and ( n12745 , n12744 , n6724 );
or ( n12746 , n12724 , n12728 , n12732 , n12736 , n12740 , n12741 , n12745 );
and ( n12747 , n12723 , n12746 );
and ( n12748 , n4027 , n3260 );
or ( n12749 , n12747 , n12748 );
and ( n12750 , n12749 , n2422 );
and ( n12751 , n4027 , n2428 );
or ( n12752 , n12750 , n12751 );
buf ( n12753 , n12752 );
buf ( n12754 , n2424 );
buf ( n12755 , n2281 );
buf ( n12756 , n2280 );
not ( n12757 , n3260 );
and ( n12758 , n4017 , n3631 );
and ( n12759 , n8819 , n5280 );
and ( n12760 , n4017 , n11909 );
or ( n12761 , n12759 , n12760 );
and ( n12762 , n12761 , n5285 );
and ( n12763 , n8830 , n5280 );
and ( n12764 , n4017 , n11909 );
or ( n12765 , n12763 , n12764 );
and ( n12766 , n12765 , n6218 );
and ( n12767 , n8841 , n5280 );
and ( n12768 , n4017 , n11909 );
or ( n12769 , n12767 , n12768 );
and ( n12770 , n12769 , n6710 );
and ( n12771 , n5514 , n5280 );
and ( n12772 , n4017 , n11909 );
or ( n12773 , n12771 , n12772 );
and ( n12774 , n12773 , n6717 );
and ( n12775 , n4015 , n6719 );
and ( n12776 , n8853 , n5280 );
and ( n12777 , n4017 , n11909 );
or ( n12778 , n12776 , n12777 );
and ( n12779 , n12778 , n6724 );
or ( n12780 , n12758 , n12762 , n12766 , n12770 , n12774 , n12775 , n12779 );
and ( n12781 , n12757 , n12780 );
and ( n12782 , n4017 , n3260 );
or ( n12783 , n12781 , n12782 );
and ( n12784 , n12783 , n2422 );
and ( n12785 , n4017 , n2428 );
nor ( n12786 , n12784 , n12785 );
buf ( n12787 , n12786 );
buf ( n12788 , n2424 );
buf ( n12789 , n2281 );
buf ( n12790 , n2280 );
not ( n12791 , n3260 );
and ( n12792 , n4007 , n3631 );
and ( n12793 , n8893 , n5280 );
and ( n12794 , n4007 , n11909 );
or ( n12795 , n12793 , n12794 );
and ( n12796 , n12795 , n5285 );
and ( n12797 , n8904 , n5280 );
and ( n12798 , n4007 , n11909 );
or ( n12799 , n12797 , n12798 );
and ( n12800 , n12799 , n6218 );
and ( n12801 , n8915 , n5280 );
and ( n12802 , n4007 , n11909 );
or ( n12803 , n12801 , n12802 );
and ( n12804 , n12803 , n6710 );
and ( n12805 , n5511 , n5280 );
and ( n12806 , n4007 , n11909 );
or ( n12807 , n12805 , n12806 );
and ( n12808 , n12807 , n6717 );
and ( n12809 , n4005 , n6719 );
and ( n12810 , n8927 , n5280 );
and ( n12811 , n4007 , n11909 );
or ( n12812 , n12810 , n12811 );
and ( n12813 , n12812 , n6724 );
or ( n12814 , n12792 , n12796 , n12800 , n12804 , n12808 , n12809 , n12813 );
and ( n12815 , n12791 , n12814 );
and ( n12816 , n4007 , n3260 );
or ( n12817 , n12815 , n12816 );
and ( n12818 , n12817 , n2422 );
and ( n12819 , n4007 , n2428 );
or ( n12820 , n12818 , n12819 );
buf ( n12821 , n12820 );
buf ( n12822 , n2424 );
buf ( n12823 , n2281 );
buf ( n12824 , n2280 );
not ( n12825 , n3260 );
and ( n12826 , n3997 , n3631 );
and ( n12827 , n8967 , n5280 );
and ( n12828 , n3997 , n11909 );
or ( n12829 , n12827 , n12828 );
and ( n12830 , n12829 , n5285 );
and ( n12831 , n8978 , n5280 );
and ( n12832 , n3997 , n11909 );
or ( n12833 , n12831 , n12832 );
and ( n12834 , n12833 , n6218 );
and ( n12835 , n8989 , n5280 );
and ( n12836 , n3997 , n11909 );
or ( n12837 , n12835 , n12836 );
and ( n12838 , n12837 , n6710 );
and ( n12839 , n5508 , n5280 );
and ( n12840 , n3997 , n11909 );
or ( n12841 , n12839 , n12840 );
and ( n12842 , n12841 , n6717 );
and ( n12843 , n3995 , n6719 );
and ( n12844 , n9001 , n5280 );
and ( n12845 , n3997 , n11909 );
or ( n12846 , n12844 , n12845 );
and ( n12847 , n12846 , n6724 );
or ( n12848 , n12826 , n12830 , n12834 , n12838 , n12842 , n12843 , n12847 );
and ( n12849 , n12825 , n12848 );
and ( n12850 , n3997 , n3260 );
or ( n12851 , n12849 , n12850 );
and ( n12852 , n12851 , n2422 );
and ( n12853 , n3997 , n2428 );
or ( n12854 , n12852 , n12853 );
buf ( n12855 , n12854 );
buf ( n12856 , n2424 );
buf ( n12857 , n2281 );
buf ( n12858 , n2280 );
not ( n12859 , n3260 );
and ( n12860 , n3987 , n3631 );
and ( n12861 , n9041 , n5280 );
and ( n12862 , n3987 , n11909 );
or ( n12863 , n12861 , n12862 );
and ( n12864 , n12863 , n5285 );
and ( n12865 , n9052 , n5280 );
and ( n12866 , n3987 , n11909 );
or ( n12867 , n12865 , n12866 );
and ( n12868 , n12867 , n6218 );
and ( n12869 , n9063 , n5280 );
and ( n12870 , n3987 , n11909 );
or ( n12871 , n12869 , n12870 );
and ( n12872 , n12871 , n6710 );
and ( n12873 , n5505 , n5280 );
and ( n12874 , n3987 , n11909 );
or ( n12875 , n12873 , n12874 );
and ( n12876 , n12875 , n6717 );
and ( n12877 , n3985 , n6719 );
and ( n12878 , n9075 , n5280 );
and ( n12879 , n3987 , n11909 );
or ( n12880 , n12878 , n12879 );
and ( n12881 , n12880 , n6724 );
or ( n12882 , n12860 , n12864 , n12868 , n12872 , n12876 , n12877 , n12881 );
and ( n12883 , n12859 , n12882 );
and ( n12884 , n3987 , n3260 );
or ( n12885 , n12883 , n12884 );
and ( n12886 , n12885 , n2422 );
and ( n12887 , n3987 , n2428 );
or ( n12888 , n12886 , n12887 );
buf ( n12889 , n12888 );
buf ( n12890 , n2424 );
buf ( n12891 , n2281 );
buf ( n12892 , n2280 );
not ( n12893 , n3260 );
and ( n12894 , n3977 , n3631 );
and ( n12895 , n10078 , n5280 );
and ( n12896 , n3977 , n11909 );
or ( n12897 , n12895 , n12896 );
and ( n12898 , n12897 , n5285 );
and ( n12899 , n10089 , n5280 );
and ( n12900 , n3977 , n11909 );
or ( n12901 , n12899 , n12900 );
and ( n12902 , n12901 , n6218 );
and ( n12903 , n10100 , n5280 );
and ( n12904 , n3977 , n11909 );
or ( n12905 , n12903 , n12904 );
and ( n12906 , n12905 , n6710 );
and ( n12907 , n5502 , n5280 );
and ( n12908 , n3977 , n11909 );
or ( n12909 , n12907 , n12908 );
and ( n12910 , n12909 , n6717 );
and ( n12911 , n3975 , n6719 );
and ( n12912 , n10111 , n5280 );
and ( n12913 , n3977 , n11909 );
or ( n12914 , n12912 , n12913 );
and ( n12915 , n12914 , n6724 );
or ( n12916 , n12894 , n12898 , n12902 , n12906 , n12910 , n12911 , n12915 );
and ( n12917 , n12893 , n12916 );
and ( n12918 , n3977 , n3260 );
or ( n12919 , n12917 , n12918 );
and ( n12920 , n12919 , n2422 );
and ( n12921 , n3977 , n2428 );
or ( n12922 , n12920 , n12921 );
buf ( n12923 , n12922 );
buf ( n12924 , n2424 );
buf ( n12925 , n2281 );
buf ( n12926 , n2280 );
not ( n12927 , n3260 );
and ( n12928 , n3813 , n3631 );
and ( n12929 , n10147 , n5280 );
and ( n12930 , n3813 , n11909 );
or ( n12931 , n12929 , n12930 );
and ( n12932 , n12931 , n5285 );
and ( n12933 , n10156 , n5280 );
and ( n12934 , n3813 , n11909 );
or ( n12935 , n12933 , n12934 );
and ( n12936 , n12935 , n6218 );
and ( n12937 , n10165 , n5280 );
and ( n12938 , n3813 , n11909 );
or ( n12939 , n12937 , n12938 );
and ( n12940 , n12939 , n6710 );
and ( n12941 , n5499 , n5280 );
and ( n12942 , n3813 , n11909 );
or ( n12943 , n12941 , n12942 );
and ( n12944 , n12943 , n6717 );
and ( n12945 , n10176 , n5280 );
and ( n12946 , n3813 , n11909 );
or ( n12947 , n12945 , n12946 );
and ( n12948 , n12947 , n6724 );
or ( n12949 , n12928 , n12932 , n12936 , n12940 , n12944 , n2424 , n12948 );
and ( n12950 , n12927 , n12949 );
and ( n12951 , n3813 , n3260 );
or ( n12952 , n12950 , n12951 );
and ( n12953 , n12952 , n2422 );
and ( n12954 , n3813 , n2428 );
or ( n12955 , n12953 , n12954 );
buf ( n12956 , n12955 );
buf ( n12957 , n2424 );
buf ( n12958 , n2281 );
buf ( n12959 , n2280 );
not ( n12960 , n3260 );
and ( n12961 , n3635 , n3631 );
and ( n12962 , n10201 , n5280 );
and ( n12963 , n3635 , n11909 );
or ( n12964 , n12962 , n12963 );
and ( n12965 , n12964 , n5285 );
and ( n12966 , n3635 , n11909 );
and ( n12967 , n12966 , n6218 );
and ( n12968 , n3635 , n11909 );
and ( n12969 , n12968 , n6710 );
and ( n12970 , n5496 , n5280 );
and ( n12971 , n3635 , n11909 );
or ( n12972 , n12970 , n12971 );
and ( n12973 , n12972 , n6717 );
and ( n12974 , n10216 , n5280 );
and ( n12975 , n3635 , n11909 );
or ( n12976 , n12974 , n12975 );
and ( n12977 , n12976 , n6724 );
or ( n12978 , n12961 , n12965 , n12967 , n12969 , n12973 , n2424 , n12977 );
and ( n12979 , n12960 , n12978 );
and ( n12980 , n3635 , n3260 );
or ( n12981 , n12979 , n12980 );
and ( n12982 , n12981 , n2422 );
and ( n12983 , n3635 , n2428 );
or ( n12984 , n12982 , n12983 );
buf ( n12985 , n12984 );
buf ( n12986 , n2424 );
buf ( n12987 , n2281 );
buf ( n12988 , n2280 );
not ( n12989 , n3066 );
not ( n12990 , n3259 );
or ( n12991 , n5285 , n3631 );
and ( n12992 , n2352 , n12991 );
xor ( n12993 , n5490 , n3789 );
not ( n12994 , n12993 );
not ( n12995 , n12994 );
and ( n12996 , n5575 , n4077 );
and ( n12997 , n5585 , n4087 );
and ( n12998 , n5595 , n4097 );
and ( n12999 , n5605 , n4107 );
and ( n13000 , n5615 , n4117 );
and ( n13001 , n5625 , n4127 );
and ( n13002 , n5635 , n4137 );
and ( n13003 , n5645 , n4147 );
and ( n13004 , n5655 , n4157 );
and ( n13005 , n5665 , n4167 );
and ( n13006 , n5675 , n4177 );
and ( n13007 , n5685 , n4187 );
and ( n13008 , n5695 , n4197 );
and ( n13009 , n5705 , n4207 );
and ( n13010 , n5715 , n4217 );
and ( n13011 , n5725 , n4227 );
and ( n13012 , n5735 , n4237 );
and ( n13013 , n5745 , n4251 );
and ( n13014 , n5755 , n3779 );
and ( n13015 , n5490 , n3789 );
and ( n13016 , n3779 , n13015 );
and ( n13017 , n5755 , n13015 );
or ( n13018 , n13014 , n13016 , n13017 );
and ( n13019 , n4251 , n13018 );
and ( n13020 , n5745 , n13018 );
or ( n13021 , n13013 , n13019 , n13020 );
and ( n13022 , n4237 , n13021 );
and ( n13023 , n5735 , n13021 );
or ( n13024 , n13012 , n13022 , n13023 );
and ( n13025 , n4227 , n13024 );
and ( n13026 , n5725 , n13024 );
or ( n13027 , n13011 , n13025 , n13026 );
and ( n13028 , n4217 , n13027 );
and ( n13029 , n5715 , n13027 );
or ( n13030 , n13010 , n13028 , n13029 );
and ( n13031 , n4207 , n13030 );
and ( n13032 , n5705 , n13030 );
or ( n13033 , n13009 , n13031 , n13032 );
and ( n13034 , n4197 , n13033 );
and ( n13035 , n5695 , n13033 );
or ( n13036 , n13008 , n13034 , n13035 );
and ( n13037 , n4187 , n13036 );
and ( n13038 , n5685 , n13036 );
or ( n13039 , n13007 , n13037 , n13038 );
and ( n13040 , n4177 , n13039 );
and ( n13041 , n5675 , n13039 );
or ( n13042 , n13006 , n13040 , n13041 );
and ( n13043 , n4167 , n13042 );
and ( n13044 , n5665 , n13042 );
or ( n13045 , n13005 , n13043 , n13044 );
and ( n13046 , n4157 , n13045 );
and ( n13047 , n5655 , n13045 );
or ( n13048 , n13004 , n13046 , n13047 );
and ( n13049 , n4147 , n13048 );
and ( n13050 , n5645 , n13048 );
or ( n13051 , n13003 , n13049 , n13050 );
and ( n13052 , n4137 , n13051 );
and ( n13053 , n5635 , n13051 );
or ( n13054 , n13002 , n13052 , n13053 );
and ( n13055 , n4127 , n13054 );
and ( n13056 , n5625 , n13054 );
or ( n13057 , n13001 , n13055 , n13056 );
and ( n13058 , n4117 , n13057 );
and ( n13059 , n5615 , n13057 );
or ( n13060 , n13000 , n13058 , n13059 );
and ( n13061 , n4107 , n13060 );
and ( n13062 , n5605 , n13060 );
or ( n13063 , n12999 , n13061 , n13062 );
and ( n13064 , n4097 , n13063 );
and ( n13065 , n5595 , n13063 );
or ( n13066 , n12998 , n13064 , n13065 );
and ( n13067 , n4087 , n13066 );
and ( n13068 , n5585 , n13066 );
or ( n13069 , n12997 , n13067 , n13068 );
and ( n13070 , n4077 , n13069 );
and ( n13071 , n5575 , n13069 );
or ( n13072 , n12996 , n13070 , n13071 );
and ( n13073 , n4067 , n13072 );
and ( n13074 , n4057 , n13073 );
and ( n13075 , n4047 , n13074 );
and ( n13076 , n4037 , n13075 );
and ( n13077 , n4027 , n13076 );
and ( n13078 , n4017 , n13077 );
and ( n13079 , n4007 , n13078 );
and ( n13080 , n3997 , n13079 );
and ( n13081 , n3987 , n13080 );
and ( n13082 , n3977 , n13081 );
and ( n13083 , n3813 , n13082 );
xor ( n13084 , n3635 , n13083 );
not ( n13085 , n13084 );
xor ( n13086 , n5755 , n3779 );
xor ( n13087 , n13086 , n13015 );
and ( n13088 , n13085 , n13087 );
not ( n13089 , n13087 );
not ( n13090 , n12993 );
xor ( n13091 , n13089 , n13090 );
and ( n13092 , n13091 , n13084 );
or ( n13093 , n13088 , n13092 );
not ( n13094 , n13093 );
not ( n13095 , n13094 );
or ( n13096 , n12995 , n13095 );
not ( n13097 , n13084 );
xor ( n13098 , n5745 , n4251 );
xor ( n13099 , n13098 , n13018 );
and ( n13100 , n13097 , n13099 );
not ( n13101 , n13099 );
and ( n13102 , n13089 , n13090 );
xor ( n13103 , n13101 , n13102 );
and ( n13104 , n13103 , n13084 );
or ( n13105 , n13100 , n13104 );
not ( n13106 , n13105 );
not ( n13107 , n13106 );
or ( n13108 , n13096 , n13107 );
not ( n13109 , n13084 );
xor ( n13110 , n5735 , n4237 );
xor ( n13111 , n13110 , n13021 );
and ( n13112 , n13109 , n13111 );
not ( n13113 , n13111 );
and ( n13114 , n13101 , n13102 );
xor ( n13115 , n13113 , n13114 );
and ( n13116 , n13115 , n13084 );
or ( n13117 , n13112 , n13116 );
not ( n13118 , n13117 );
not ( n13119 , n13118 );
or ( n13120 , n13108 , n13119 );
not ( n13121 , n13084 );
xor ( n13122 , n5725 , n4227 );
xor ( n13123 , n13122 , n13024 );
and ( n13124 , n13121 , n13123 );
not ( n13125 , n13123 );
and ( n13126 , n13113 , n13114 );
xor ( n13127 , n13125 , n13126 );
and ( n13128 , n13127 , n13084 );
or ( n13129 , n13124 , n13128 );
not ( n13130 , n13129 );
not ( n13131 , n13130 );
or ( n13132 , n13120 , n13131 );
not ( n13133 , n13084 );
xor ( n13134 , n5715 , n4217 );
xor ( n13135 , n13134 , n13027 );
and ( n13136 , n13133 , n13135 );
not ( n13137 , n13135 );
and ( n13138 , n13125 , n13126 );
xor ( n13139 , n13137 , n13138 );
and ( n13140 , n13139 , n13084 );
or ( n13141 , n13136 , n13140 );
not ( n13142 , n13141 );
not ( n13143 , n13142 );
or ( n13144 , n13132 , n13143 );
not ( n13145 , n13084 );
xor ( n13146 , n5705 , n4207 );
xor ( n13147 , n13146 , n13030 );
and ( n13148 , n13145 , n13147 );
not ( n13149 , n13147 );
and ( n13150 , n13137 , n13138 );
xor ( n13151 , n13149 , n13150 );
and ( n13152 , n13151 , n13084 );
or ( n13153 , n13148 , n13152 );
not ( n13154 , n13153 );
not ( n13155 , n13154 );
or ( n13156 , n13144 , n13155 );
not ( n13157 , n13084 );
xor ( n13158 , n5695 , n4197 );
xor ( n13159 , n13158 , n13033 );
and ( n13160 , n13157 , n13159 );
not ( n13161 , n13159 );
and ( n13162 , n13149 , n13150 );
xor ( n13163 , n13161 , n13162 );
and ( n13164 , n13163 , n13084 );
or ( n13165 , n13160 , n13164 );
not ( n13166 , n13165 );
not ( n13167 , n13166 );
or ( n13168 , n13156 , n13167 );
not ( n13169 , n13084 );
xor ( n13170 , n5685 , n4187 );
xor ( n13171 , n13170 , n13036 );
and ( n13172 , n13169 , n13171 );
not ( n13173 , n13171 );
and ( n13174 , n13161 , n13162 );
xor ( n13175 , n13173 , n13174 );
and ( n13176 , n13175 , n13084 );
or ( n13177 , n13172 , n13176 );
not ( n13178 , n13177 );
not ( n13179 , n13178 );
or ( n13180 , n13168 , n13179 );
not ( n13181 , n13084 );
xor ( n13182 , n5675 , n4177 );
xor ( n13183 , n13182 , n13039 );
and ( n13184 , n13181 , n13183 );
not ( n13185 , n13183 );
and ( n13186 , n13173 , n13174 );
xor ( n13187 , n13185 , n13186 );
and ( n13188 , n13187 , n13084 );
or ( n13189 , n13184 , n13188 );
not ( n13190 , n13189 );
not ( n13191 , n13190 );
or ( n13192 , n13180 , n13191 );
not ( n13193 , n13084 );
xor ( n13194 , n5665 , n4167 );
xor ( n13195 , n13194 , n13042 );
and ( n13196 , n13193 , n13195 );
not ( n13197 , n13195 );
and ( n13198 , n13185 , n13186 );
xor ( n13199 , n13197 , n13198 );
and ( n13200 , n13199 , n13084 );
or ( n13201 , n13196 , n13200 );
not ( n13202 , n13201 );
not ( n13203 , n13202 );
or ( n13204 , n13192 , n13203 );
not ( n13205 , n13084 );
xor ( n13206 , n5655 , n4157 );
xor ( n13207 , n13206 , n13045 );
and ( n13208 , n13205 , n13207 );
not ( n13209 , n13207 );
and ( n13210 , n13197 , n13198 );
xor ( n13211 , n13209 , n13210 );
and ( n13212 , n13211 , n13084 );
or ( n13213 , n13208 , n13212 );
not ( n13214 , n13213 );
not ( n13215 , n13214 );
or ( n13216 , n13204 , n13215 );
not ( n13217 , n13084 );
xor ( n13218 , n5645 , n4147 );
xor ( n13219 , n13218 , n13048 );
and ( n13220 , n13217 , n13219 );
not ( n13221 , n13219 );
and ( n13222 , n13209 , n13210 );
xor ( n13223 , n13221 , n13222 );
and ( n13224 , n13223 , n13084 );
or ( n13225 , n13220 , n13224 );
not ( n13226 , n13225 );
not ( n13227 , n13226 );
or ( n13228 , n13216 , n13227 );
not ( n13229 , n13084 );
xor ( n13230 , n5635 , n4137 );
xor ( n13231 , n13230 , n13051 );
and ( n13232 , n13229 , n13231 );
not ( n13233 , n13231 );
and ( n13234 , n13221 , n13222 );
xor ( n13235 , n13233 , n13234 );
and ( n13236 , n13235 , n13084 );
or ( n13237 , n13232 , n13236 );
not ( n13238 , n13237 );
not ( n13239 , n13238 );
or ( n13240 , n13228 , n13239 );
not ( n13241 , n13084 );
xor ( n13242 , n5625 , n4127 );
xor ( n13243 , n13242 , n13054 );
and ( n13244 , n13241 , n13243 );
not ( n13245 , n13243 );
and ( n13246 , n13233 , n13234 );
xor ( n13247 , n13245 , n13246 );
and ( n13248 , n13247 , n13084 );
or ( n13249 , n13244 , n13248 );
not ( n13250 , n13249 );
not ( n13251 , n13250 );
xor ( n13252 , n13240 , n13251 );
not ( n13253 , n13084 );
xor ( n13254 , n5615 , n4117 );
xor ( n13255 , n13254 , n13057 );
and ( n13256 , n13253 , n13255 );
not ( n13257 , n13255 );
and ( n13258 , n13245 , n13246 );
xor ( n13259 , n13257 , n13258 );
and ( n13260 , n13259 , n13084 );
or ( n13261 , n13256 , n13260 );
not ( n13262 , n13261 );
not ( n13263 , n13262 );
or ( n13264 , n13252 , n13263 );
not ( n13265 , n13084 );
xor ( n13266 , n5605 , n4107 );
xor ( n13267 , n13266 , n13060 );
and ( n13268 , n13265 , n13267 );
not ( n13269 , n13267 );
and ( n13270 , n13257 , n13258 );
xor ( n13271 , n13269 , n13270 );
and ( n13272 , n13271 , n13084 );
or ( n13273 , n13268 , n13272 );
not ( n13274 , n13273 );
not ( n13275 , n13274 );
or ( n13276 , n13264 , n13275 );
not ( n13277 , n13084 );
xor ( n13278 , n5595 , n4097 );
xor ( n13279 , n13278 , n13063 );
and ( n13280 , n13277 , n13279 );
not ( n13281 , n13279 );
and ( n13282 , n13269 , n13270 );
xor ( n13283 , n13281 , n13282 );
and ( n13284 , n13283 , n13084 );
or ( n13285 , n13280 , n13284 );
not ( n13286 , n13285 );
not ( n13287 , n13286 );
or ( n13288 , n13276 , n13287 );
not ( n13289 , n13084 );
xor ( n13290 , n5585 , n4087 );
xor ( n13291 , n13290 , n13066 );
and ( n13292 , n13289 , n13291 );
not ( n13293 , n13291 );
and ( n13294 , n13281 , n13282 );
xor ( n13295 , n13293 , n13294 );
and ( n13296 , n13295 , n13084 );
or ( n13297 , n13292 , n13296 );
not ( n13298 , n13297 );
not ( n13299 , n13298 );
or ( n13300 , n13288 , n13299 );
not ( n13301 , n13084 );
xor ( n13302 , n5575 , n4077 );
xor ( n13303 , n13302 , n13069 );
and ( n13304 , n13301 , n13303 );
not ( n13305 , n13303 );
and ( n13306 , n13293 , n13294 );
xor ( n13307 , n13305 , n13306 );
and ( n13308 , n13307 , n13084 );
or ( n13309 , n13304 , n13308 );
not ( n13310 , n13309 );
not ( n13311 , n13310 );
or ( n13312 , n13300 , n13311 );
and ( n13313 , n13312 , n13084 );
not ( n13314 , n13313 );
and ( n13315 , n13314 , n12995 );
xor ( n13316 , n12995 , n13084 );
xor ( n13317 , n13316 , n13084 );
and ( n13318 , n13317 , n13313 );
or ( n13319 , n13315 , n13318 );
and ( n13320 , n13319 , n5289 );
xor ( n13321 , n5490 , n3791 );
not ( n13322 , n13321 );
not ( n13323 , n13322 );
and ( n13324 , n5575 , n4079 );
and ( n13325 , n5585 , n4089 );
and ( n13326 , n5595 , n4099 );
and ( n13327 , n5605 , n4109 );
and ( n13328 , n5615 , n4119 );
and ( n13329 , n5625 , n4129 );
and ( n13330 , n5635 , n4139 );
and ( n13331 , n5645 , n4149 );
and ( n13332 , n5655 , n4159 );
and ( n13333 , n5665 , n4169 );
and ( n13334 , n5675 , n4179 );
and ( n13335 , n5685 , n4189 );
and ( n13336 , n5695 , n4199 );
and ( n13337 , n5705 , n4209 );
and ( n13338 , n5715 , n4219 );
and ( n13339 , n5725 , n4229 );
and ( n13340 , n5735 , n4239 );
and ( n13341 , n5745 , n4253 );
and ( n13342 , n5755 , n3781 );
and ( n13343 , n5490 , n3791 );
and ( n13344 , n3781 , n13343 );
and ( n13345 , n5755 , n13343 );
or ( n13346 , n13342 , n13344 , n13345 );
and ( n13347 , n4253 , n13346 );
and ( n13348 , n5745 , n13346 );
or ( n13349 , n13341 , n13347 , n13348 );
and ( n13350 , n4239 , n13349 );
and ( n13351 , n5735 , n13349 );
or ( n13352 , n13340 , n13350 , n13351 );
and ( n13353 , n4229 , n13352 );
and ( n13354 , n5725 , n13352 );
or ( n13355 , n13339 , n13353 , n13354 );
and ( n13356 , n4219 , n13355 );
and ( n13357 , n5715 , n13355 );
or ( n13358 , n13338 , n13356 , n13357 );
and ( n13359 , n4209 , n13358 );
and ( n13360 , n5705 , n13358 );
or ( n13361 , n13337 , n13359 , n13360 );
and ( n13362 , n4199 , n13361 );
and ( n13363 , n5695 , n13361 );
or ( n13364 , n13336 , n13362 , n13363 );
and ( n13365 , n4189 , n13364 );
and ( n13366 , n5685 , n13364 );
or ( n13367 , n13335 , n13365 , n13366 );
and ( n13368 , n4179 , n13367 );
and ( n13369 , n5675 , n13367 );
or ( n13370 , n13334 , n13368 , n13369 );
and ( n13371 , n4169 , n13370 );
and ( n13372 , n5665 , n13370 );
or ( n13373 , n13333 , n13371 , n13372 );
and ( n13374 , n4159 , n13373 );
and ( n13375 , n5655 , n13373 );
or ( n13376 , n13332 , n13374 , n13375 );
and ( n13377 , n4149 , n13376 );
and ( n13378 , n5645 , n13376 );
or ( n13379 , n13331 , n13377 , n13378 );
and ( n13380 , n4139 , n13379 );
and ( n13381 , n5635 , n13379 );
or ( n13382 , n13330 , n13380 , n13381 );
and ( n13383 , n4129 , n13382 );
and ( n13384 , n5625 , n13382 );
or ( n13385 , n13329 , n13383 , n13384 );
and ( n13386 , n4119 , n13385 );
and ( n13387 , n5615 , n13385 );
or ( n13388 , n13328 , n13386 , n13387 );
and ( n13389 , n4109 , n13388 );
and ( n13390 , n5605 , n13388 );
or ( n13391 , n13327 , n13389 , n13390 );
and ( n13392 , n4099 , n13391 );
and ( n13393 , n5595 , n13391 );
or ( n13394 , n13326 , n13392 , n13393 );
and ( n13395 , n4089 , n13394 );
and ( n13396 , n5585 , n13394 );
or ( n13397 , n13325 , n13395 , n13396 );
and ( n13398 , n4079 , n13397 );
and ( n13399 , n5575 , n13397 );
or ( n13400 , n13324 , n13398 , n13399 );
and ( n13401 , n4069 , n13400 );
and ( n13402 , n4059 , n13401 );
and ( n13403 , n4049 , n13402 );
and ( n13404 , n4039 , n13403 );
and ( n13405 , n4029 , n13404 );
and ( n13406 , n4019 , n13405 );
and ( n13407 , n4009 , n13406 );
and ( n13408 , n3999 , n13407 );
and ( n13409 , n3989 , n13408 );
and ( n13410 , n3979 , n13409 );
and ( n13411 , n3815 , n13410 );
xor ( n13412 , n3764 , n13411 );
not ( n13413 , n13412 );
xor ( n13414 , n5755 , n3781 );
xor ( n13415 , n13414 , n13343 );
and ( n13416 , n13413 , n13415 );
not ( n13417 , n13415 );
not ( n13418 , n13321 );
xor ( n13419 , n13417 , n13418 );
and ( n13420 , n13419 , n13412 );
or ( n13421 , n13416 , n13420 );
not ( n13422 , n13421 );
not ( n13423 , n13422 );
or ( n13424 , n13323 , n13423 );
not ( n13425 , n13412 );
xor ( n13426 , n5745 , n4253 );
xor ( n13427 , n13426 , n13346 );
and ( n13428 , n13425 , n13427 );
not ( n13429 , n13427 );
and ( n13430 , n13417 , n13418 );
xor ( n13431 , n13429 , n13430 );
and ( n13432 , n13431 , n13412 );
or ( n13433 , n13428 , n13432 );
not ( n13434 , n13433 );
not ( n13435 , n13434 );
or ( n13436 , n13424 , n13435 );
not ( n13437 , n13412 );
xor ( n13438 , n5735 , n4239 );
xor ( n13439 , n13438 , n13349 );
and ( n13440 , n13437 , n13439 );
not ( n13441 , n13439 );
and ( n13442 , n13429 , n13430 );
xor ( n13443 , n13441 , n13442 );
and ( n13444 , n13443 , n13412 );
or ( n13445 , n13440 , n13444 );
not ( n13446 , n13445 );
not ( n13447 , n13446 );
or ( n13448 , n13436 , n13447 );
not ( n13449 , n13412 );
xor ( n13450 , n5725 , n4229 );
xor ( n13451 , n13450 , n13352 );
and ( n13452 , n13449 , n13451 );
not ( n13453 , n13451 );
and ( n13454 , n13441 , n13442 );
xor ( n13455 , n13453 , n13454 );
and ( n13456 , n13455 , n13412 );
or ( n13457 , n13452 , n13456 );
not ( n13458 , n13457 );
not ( n13459 , n13458 );
or ( n13460 , n13448 , n13459 );
not ( n13461 , n13412 );
xor ( n13462 , n5715 , n4219 );
xor ( n13463 , n13462 , n13355 );
and ( n13464 , n13461 , n13463 );
not ( n13465 , n13463 );
and ( n13466 , n13453 , n13454 );
xor ( n13467 , n13465 , n13466 );
and ( n13468 , n13467 , n13412 );
or ( n13469 , n13464 , n13468 );
not ( n13470 , n13469 );
not ( n13471 , n13470 );
or ( n13472 , n13460 , n13471 );
not ( n13473 , n13412 );
xor ( n13474 , n5705 , n4209 );
xor ( n13475 , n13474 , n13358 );
and ( n13476 , n13473 , n13475 );
not ( n13477 , n13475 );
and ( n13478 , n13465 , n13466 );
xor ( n13479 , n13477 , n13478 );
and ( n13480 , n13479 , n13412 );
or ( n13481 , n13476 , n13480 );
not ( n13482 , n13481 );
not ( n13483 , n13482 );
or ( n13484 , n13472 , n13483 );
not ( n13485 , n13412 );
xor ( n13486 , n5695 , n4199 );
xor ( n13487 , n13486 , n13361 );
and ( n13488 , n13485 , n13487 );
not ( n13489 , n13487 );
and ( n13490 , n13477 , n13478 );
xor ( n13491 , n13489 , n13490 );
and ( n13492 , n13491 , n13412 );
or ( n13493 , n13488 , n13492 );
not ( n13494 , n13493 );
not ( n13495 , n13494 );
or ( n13496 , n13484 , n13495 );
not ( n13497 , n13412 );
xor ( n13498 , n5685 , n4189 );
xor ( n13499 , n13498 , n13364 );
and ( n13500 , n13497 , n13499 );
not ( n13501 , n13499 );
and ( n13502 , n13489 , n13490 );
xor ( n13503 , n13501 , n13502 );
and ( n13504 , n13503 , n13412 );
or ( n13505 , n13500 , n13504 );
not ( n13506 , n13505 );
not ( n13507 , n13506 );
or ( n13508 , n13496 , n13507 );
not ( n13509 , n13412 );
xor ( n13510 , n5675 , n4179 );
xor ( n13511 , n13510 , n13367 );
and ( n13512 , n13509 , n13511 );
not ( n13513 , n13511 );
and ( n13514 , n13501 , n13502 );
xor ( n13515 , n13513 , n13514 );
and ( n13516 , n13515 , n13412 );
or ( n13517 , n13512 , n13516 );
not ( n13518 , n13517 );
not ( n13519 , n13518 );
or ( n13520 , n13508 , n13519 );
not ( n13521 , n13412 );
xor ( n13522 , n5665 , n4169 );
xor ( n13523 , n13522 , n13370 );
and ( n13524 , n13521 , n13523 );
not ( n13525 , n13523 );
and ( n13526 , n13513 , n13514 );
xor ( n13527 , n13525 , n13526 );
and ( n13528 , n13527 , n13412 );
or ( n13529 , n13524 , n13528 );
not ( n13530 , n13529 );
not ( n13531 , n13530 );
or ( n13532 , n13520 , n13531 );
not ( n13533 , n13412 );
xor ( n13534 , n5655 , n4159 );
xor ( n13535 , n13534 , n13373 );
and ( n13536 , n13533 , n13535 );
not ( n13537 , n13535 );
and ( n13538 , n13525 , n13526 );
xor ( n13539 , n13537 , n13538 );
and ( n13540 , n13539 , n13412 );
or ( n13541 , n13536 , n13540 );
not ( n13542 , n13541 );
not ( n13543 , n13542 );
or ( n13544 , n13532 , n13543 );
not ( n13545 , n13412 );
xor ( n13546 , n5645 , n4149 );
xor ( n13547 , n13546 , n13376 );
and ( n13548 , n13545 , n13547 );
not ( n13549 , n13547 );
and ( n13550 , n13537 , n13538 );
xor ( n13551 , n13549 , n13550 );
and ( n13552 , n13551 , n13412 );
or ( n13553 , n13548 , n13552 );
not ( n13554 , n13553 );
not ( n13555 , n13554 );
or ( n13556 , n13544 , n13555 );
not ( n13557 , n13412 );
xor ( n13558 , n5635 , n4139 );
xor ( n13559 , n13558 , n13379 );
and ( n13560 , n13557 , n13559 );
not ( n13561 , n13559 );
and ( n13562 , n13549 , n13550 );
xor ( n13563 , n13561 , n13562 );
and ( n13564 , n13563 , n13412 );
or ( n13565 , n13560 , n13564 );
not ( n13566 , n13565 );
not ( n13567 , n13566 );
or ( n13568 , n13556 , n13567 );
not ( n13569 , n13412 );
xor ( n13570 , n5625 , n4129 );
xor ( n13571 , n13570 , n13382 );
and ( n13572 , n13569 , n13571 );
not ( n13573 , n13571 );
and ( n13574 , n13561 , n13562 );
xor ( n13575 , n13573 , n13574 );
and ( n13576 , n13575 , n13412 );
or ( n13577 , n13572 , n13576 );
not ( n13578 , n13577 );
not ( n13579 , n13578 );
or ( n13580 , n13568 , n13579 );
not ( n13581 , n13412 );
xor ( n13582 , n5615 , n4119 );
xor ( n13583 , n13582 , n13385 );
and ( n13584 , n13581 , n13583 );
not ( n13585 , n13583 );
and ( n13586 , n13573 , n13574 );
xor ( n13587 , n13585 , n13586 );
and ( n13588 , n13587 , n13412 );
or ( n13589 , n13584 , n13588 );
not ( n13590 , n13589 );
not ( n13591 , n13590 );
or ( n13592 , n13580 , n13591 );
not ( n13593 , n13412 );
xor ( n13594 , n5605 , n4109 );
xor ( n13595 , n13594 , n13388 );
and ( n13596 , n13593 , n13595 );
not ( n13597 , n13595 );
and ( n13598 , n13585 , n13586 );
xor ( n13599 , n13597 , n13598 );
and ( n13600 , n13599 , n13412 );
or ( n13601 , n13596 , n13600 );
not ( n13602 , n13601 );
not ( n13603 , n13602 );
or ( n13604 , n13592 , n13603 );
not ( n13605 , n13412 );
xor ( n13606 , n5595 , n4099 );
xor ( n13607 , n13606 , n13391 );
and ( n13608 , n13605 , n13607 );
not ( n13609 , n13607 );
and ( n13610 , n13597 , n13598 );
xor ( n13611 , n13609 , n13610 );
and ( n13612 , n13611 , n13412 );
or ( n13613 , n13608 , n13612 );
not ( n13614 , n13613 );
not ( n13615 , n13614 );
or ( n13616 , n13604 , n13615 );
not ( n13617 , n13412 );
xor ( n13618 , n5585 , n4089 );
xor ( n13619 , n13618 , n13394 );
and ( n13620 , n13617 , n13619 );
not ( n13621 , n13619 );
and ( n13622 , n13609 , n13610 );
xor ( n13623 , n13621 , n13622 );
and ( n13624 , n13623 , n13412 );
or ( n13625 , n13620 , n13624 );
not ( n13626 , n13625 );
not ( n13627 , n13626 );
or ( n13628 , n13616 , n13627 );
not ( n13629 , n13412 );
xor ( n13630 , n5575 , n4079 );
xor ( n13631 , n13630 , n13397 );
and ( n13632 , n13629 , n13631 );
not ( n13633 , n13631 );
and ( n13634 , n13621 , n13622 );
xor ( n13635 , n13633 , n13634 );
and ( n13636 , n13635 , n13412 );
or ( n13637 , n13632 , n13636 );
not ( n13638 , n13637 );
not ( n13639 , n13638 );
or ( n13640 , n13628 , n13639 );
and ( n13641 , n13640 , n13412 );
not ( n13642 , n13641 );
and ( n13643 , n13642 , n13323 );
xor ( n13644 , n13323 , n13412 );
xor ( n13645 , n13644 , n13412 );
and ( n13646 , n13645 , n13641 );
or ( n13647 , n13643 , n13646 );
and ( n13648 , n13647 , n5287 );
and ( n13649 , n5490 , n5152 );
and ( n13650 , n2352 , n5154 );
or ( n13651 , n13320 , n13648 , n13649 , n13650 );
or ( n13652 , n6724 , n6719 );
or ( n13653 , n13652 , n6715 );
or ( n13654 , n13653 , n6716 );
or ( n13655 , n13654 , n6704 );
or ( n13656 , n13655 , n6705 );
or ( n13657 , n13656 , n6212 );
or ( n13658 , n13657 , n6213 );
or ( n13659 , n13658 , n6707 );
or ( n13660 , n13659 , n6215 );
or ( n13661 , n13660 , n6709 );
or ( n13662 , n13661 , n6217 );
and ( n13663 , n13651 , n13662 );
or ( n13664 , n12992 , n13663 );
and ( n13665 , n12990 , n13664 );
and ( n13666 , n2424 , n3259 );
or ( n13667 , n13665 , n13666 );
and ( n13668 , n12989 , n13667 );
and ( n13669 , n13651 , n3066 );
or ( n13670 , n13668 , n13669 );
and ( n13671 , n13670 , n2422 );
not ( n13672 , n3356 );
not ( n13673 , n13672 );
buf ( n13674 , n13673 );
and ( n13675 , n13674 , n2428 );
or ( n13676 , n13671 , n13675 );
buf ( n13677 , n13676 );
buf ( n13678 , n2424 );
buf ( n13679 , n2281 );
buf ( n13680 , n2280 );
not ( n13681 , n3066 );
not ( n13682 , n3259 );
and ( n13683 , n2350 , n12991 );
not ( n13684 , n13313 );
and ( n13685 , n13684 , n13095 );
xor ( n13686 , n13095 , n13084 );
and ( n13687 , n13316 , n13084 );
xor ( n13688 , n13686 , n13687 );
and ( n13689 , n13688 , n13313 );
or ( n13690 , n13685 , n13689 );
and ( n13691 , n13690 , n5289 );
not ( n13692 , n13641 );
and ( n13693 , n13692 , n13423 );
xor ( n13694 , n13423 , n13412 );
and ( n13695 , n13644 , n13412 );
xor ( n13696 , n13694 , n13695 );
and ( n13697 , n13696 , n13641 );
or ( n13698 , n13693 , n13697 );
and ( n13699 , n13698 , n5287 );
and ( n13700 , n5755 , n5152 );
and ( n13701 , n2350 , n5154 );
or ( n13702 , n13691 , n13699 , n13700 , n13701 );
and ( n13703 , n13702 , n13662 );
or ( n13704 , n13683 , n13703 );
and ( n13705 , n13682 , n13704 );
and ( n13706 , n2424 , n3259 );
or ( n13707 , n13705 , n13706 );
and ( n13708 , n13681 , n13707 );
and ( n13709 , n13702 , n3066 );
or ( n13710 , n13708 , n13709 );
and ( n13711 , n13710 , n2422 );
buf ( n13712 , n3772 );
not ( n13713 , n13712 );
not ( n13714 , n13713 );
buf ( n13715 , n13714 );
and ( n13716 , n13715 , n2428 );
or ( n13717 , n13711 , n13716 );
buf ( n13718 , n13717 );
buf ( n13719 , n2424 );
buf ( n13720 , n2281 );
buf ( n13721 , n2280 );
not ( n13722 , n3066 );
not ( n13723 , n3259 );
and ( n13724 , n2348 , n12991 );
not ( n13725 , n13313 );
and ( n13726 , n13725 , n13107 );
xor ( n13727 , n13107 , n13084 );
and ( n13728 , n13686 , n13687 );
xor ( n13729 , n13727 , n13728 );
and ( n13730 , n13729 , n13313 );
or ( n13731 , n13726 , n13730 );
and ( n13732 , n13731 , n5289 );
not ( n13733 , n13641 );
and ( n13734 , n13733 , n13435 );
xor ( n13735 , n13435 , n13412 );
and ( n13736 , n13694 , n13695 );
xor ( n13737 , n13735 , n13736 );
and ( n13738 , n13737 , n13641 );
or ( n13739 , n13734 , n13738 );
and ( n13740 , n13739 , n5287 );
and ( n13741 , n5745 , n5152 );
and ( n13742 , n2348 , n5154 );
or ( n13743 , n13732 , n13740 , n13741 , n13742 );
and ( n13744 , n13743 , n13662 );
or ( n13745 , n13724 , n13744 );
and ( n13746 , n13723 , n13745 );
not ( n13747 , n3789 );
not ( n13748 , n13747 );
not ( n13749 , n3635 );
and ( n13750 , n13749 , n3779 );
not ( n13751 , n3779 );
not ( n13752 , n3789 );
xor ( n13753 , n13751 , n13752 );
and ( n13754 , n13753 , n3635 );
or ( n13755 , n13750 , n13754 );
not ( n13756 , n13755 );
not ( n13757 , n13756 );
or ( n13758 , n13748 , n13757 );
not ( n13759 , n3635 );
and ( n13760 , n13759 , n4251 );
not ( n13761 , n4251 );
and ( n13762 , n13751 , n13752 );
xor ( n13763 , n13761 , n13762 );
and ( n13764 , n13763 , n3635 );
or ( n13765 , n13760 , n13764 );
not ( n13766 , n13765 );
not ( n13767 , n13766 );
or ( n13768 , n13758 , n13767 );
not ( n13769 , n3635 );
and ( n13770 , n13769 , n4237 );
not ( n13771 , n4237 );
and ( n13772 , n13761 , n13762 );
xor ( n13773 , n13771 , n13772 );
and ( n13774 , n13773 , n3635 );
or ( n13775 , n13770 , n13774 );
not ( n13776 , n13775 );
not ( n13777 , n13776 );
or ( n13778 , n13768 , n13777 );
not ( n13779 , n3635 );
and ( n13780 , n13779 , n4227 );
not ( n13781 , n4227 );
and ( n13782 , n13771 , n13772 );
xor ( n13783 , n13781 , n13782 );
and ( n13784 , n13783 , n3635 );
or ( n13785 , n13780 , n13784 );
not ( n13786 , n13785 );
not ( n13787 , n13786 );
or ( n13788 , n13778 , n13787 );
not ( n13789 , n3635 );
and ( n13790 , n13789 , n4217 );
not ( n13791 , n4217 );
and ( n13792 , n13781 , n13782 );
xor ( n13793 , n13791 , n13792 );
and ( n13794 , n13793 , n3635 );
or ( n13795 , n13790 , n13794 );
not ( n13796 , n13795 );
not ( n13797 , n13796 );
or ( n13798 , n13788 , n13797 );
not ( n13799 , n3635 );
and ( n13800 , n13799 , n4207 );
not ( n13801 , n4207 );
and ( n13802 , n13791 , n13792 );
xor ( n13803 , n13801 , n13802 );
and ( n13804 , n13803 , n3635 );
or ( n13805 , n13800 , n13804 );
not ( n13806 , n13805 );
not ( n13807 , n13806 );
or ( n13808 , n13798 , n13807 );
not ( n13809 , n3635 );
and ( n13810 , n13809 , n4197 );
not ( n13811 , n4197 );
and ( n13812 , n13801 , n13802 );
xor ( n13813 , n13811 , n13812 );
and ( n13814 , n13813 , n3635 );
or ( n13815 , n13810 , n13814 );
not ( n13816 , n13815 );
not ( n13817 , n13816 );
or ( n13818 , n13808 , n13817 );
not ( n13819 , n3635 );
and ( n13820 , n13819 , n4187 );
not ( n13821 , n4187 );
and ( n13822 , n13811 , n13812 );
xor ( n13823 , n13821 , n13822 );
and ( n13824 , n13823 , n3635 );
or ( n13825 , n13820 , n13824 );
not ( n13826 , n13825 );
not ( n13827 , n13826 );
or ( n13828 , n13818 , n13827 );
not ( n13829 , n3635 );
and ( n13830 , n13829 , n4177 );
not ( n13831 , n4177 );
and ( n13832 , n13821 , n13822 );
xor ( n13833 , n13831 , n13832 );
and ( n13834 , n13833 , n3635 );
or ( n13835 , n13830 , n13834 );
not ( n13836 , n13835 );
not ( n13837 , n13836 );
or ( n13838 , n13828 , n13837 );
not ( n13839 , n3635 );
and ( n13840 , n13839 , n4167 );
not ( n13841 , n4167 );
and ( n13842 , n13831 , n13832 );
xor ( n13843 , n13841 , n13842 );
and ( n13844 , n13843 , n3635 );
or ( n13845 , n13840 , n13844 );
not ( n13846 , n13845 );
not ( n13847 , n13846 );
or ( n13848 , n13838 , n13847 );
not ( n13849 , n3635 );
and ( n13850 , n13849 , n4157 );
not ( n13851 , n4157 );
and ( n13852 , n13841 , n13842 );
xor ( n13853 , n13851 , n13852 );
and ( n13854 , n13853 , n3635 );
or ( n13855 , n13850 , n13854 );
not ( n13856 , n13855 );
not ( n13857 , n13856 );
or ( n13858 , n13848 , n13857 );
not ( n13859 , n3635 );
and ( n13860 , n13859 , n4147 );
not ( n13861 , n4147 );
and ( n13862 , n13851 , n13852 );
xor ( n13863 , n13861 , n13862 );
and ( n13864 , n13863 , n3635 );
or ( n13865 , n13860 , n13864 );
not ( n13866 , n13865 );
not ( n13867 , n13866 );
or ( n13868 , n13858 , n13867 );
not ( n13869 , n3635 );
and ( n13870 , n13869 , n4137 );
not ( n13871 , n4137 );
and ( n13872 , n13861 , n13862 );
xor ( n13873 , n13871 , n13872 );
and ( n13874 , n13873 , n3635 );
or ( n13875 , n13870 , n13874 );
not ( n13876 , n13875 );
not ( n13877 , n13876 );
or ( n13878 , n13868 , n13877 );
not ( n13879 , n3635 );
and ( n13880 , n13879 , n4127 );
not ( n13881 , n4127 );
and ( n13882 , n13871 , n13872 );
xor ( n13883 , n13881 , n13882 );
and ( n13884 , n13883 , n3635 );
or ( n13885 , n13880 , n13884 );
not ( n13886 , n13885 );
not ( n13887 , n13886 );
or ( n13888 , n13878 , n13887 );
not ( n13889 , n3635 );
and ( n13890 , n13889 , n4117 );
not ( n13891 , n4117 );
and ( n13892 , n13881 , n13882 );
xor ( n13893 , n13891 , n13892 );
and ( n13894 , n13893 , n3635 );
or ( n13895 , n13890 , n13894 );
not ( n13896 , n13895 );
not ( n13897 , n13896 );
or ( n13898 , n13888 , n13897 );
not ( n13899 , n3635 );
and ( n13900 , n13899 , n4107 );
not ( n13901 , n4107 );
and ( n13902 , n13891 , n13892 );
xor ( n13903 , n13901 , n13902 );
and ( n13904 , n13903 , n3635 );
or ( n13905 , n13900 , n13904 );
not ( n13906 , n13905 );
not ( n13907 , n13906 );
or ( n13908 , n13898 , n13907 );
not ( n13909 , n3635 );
and ( n13910 , n13909 , n4097 );
not ( n13911 , n4097 );
and ( n13912 , n13901 , n13902 );
xor ( n13913 , n13911 , n13912 );
and ( n13914 , n13913 , n3635 );
or ( n13915 , n13910 , n13914 );
not ( n13916 , n13915 );
not ( n13917 , n13916 );
or ( n13918 , n13908 , n13917 );
not ( n13919 , n3635 );
and ( n13920 , n13919 , n4087 );
not ( n13921 , n4087 );
and ( n13922 , n13911 , n13912 );
xor ( n13923 , n13921 , n13922 );
and ( n13924 , n13923 , n3635 );
or ( n13925 , n13920 , n13924 );
not ( n13926 , n13925 );
not ( n13927 , n13926 );
or ( n13928 , n13918 , n13927 );
not ( n13929 , n3635 );
and ( n13930 , n13929 , n4077 );
not ( n13931 , n4077 );
and ( n13932 , n13921 , n13922 );
xor ( n13933 , n13931 , n13932 );
and ( n13934 , n13933 , n3635 );
or ( n13935 , n13930 , n13934 );
not ( n13936 , n13935 );
not ( n13937 , n13936 );
or ( n13938 , n13928 , n13937 );
and ( n13939 , n13938 , n3635 );
not ( n13940 , n13939 );
and ( n13941 , n13940 , n13748 );
xor ( n13942 , n13748 , n3635 );
xor ( n13943 , n13942 , n3635 );
and ( n13944 , n13943 , n13939 );
or ( n13945 , n13941 , n13944 );
not ( n13946 , n5490 );
not ( n13947 , n13946 );
xor ( n13948 , n13945 , n13947 );
and ( n13949 , n13948 , n5289 );
not ( n13950 , n3791 );
not ( n13951 , n13950 );
not ( n13952 , n3764 );
and ( n13953 , n13952 , n3781 );
not ( n13954 , n3781 );
not ( n13955 , n3791 );
xor ( n13956 , n13954 , n13955 );
and ( n13957 , n13956 , n3764 );
or ( n13958 , n13953 , n13957 );
not ( n13959 , n13958 );
not ( n13960 , n13959 );
or ( n13961 , n13951 , n13960 );
not ( n13962 , n3764 );
and ( n13963 , n13962 , n4253 );
not ( n13964 , n4253 );
and ( n13965 , n13954 , n13955 );
xor ( n13966 , n13964 , n13965 );
and ( n13967 , n13966 , n3764 );
or ( n13968 , n13963 , n13967 );
not ( n13969 , n13968 );
not ( n13970 , n13969 );
or ( n13971 , n13961 , n13970 );
not ( n13972 , n3764 );
and ( n13973 , n13972 , n4239 );
not ( n13974 , n4239 );
and ( n13975 , n13964 , n13965 );
xor ( n13976 , n13974 , n13975 );
and ( n13977 , n13976 , n3764 );
or ( n13978 , n13973 , n13977 );
not ( n13979 , n13978 );
not ( n13980 , n13979 );
or ( n13981 , n13971 , n13980 );
not ( n13982 , n3764 );
and ( n13983 , n13982 , n4229 );
not ( n13984 , n4229 );
and ( n13985 , n13974 , n13975 );
xor ( n13986 , n13984 , n13985 );
and ( n13987 , n13986 , n3764 );
or ( n13988 , n13983 , n13987 );
not ( n13989 , n13988 );
not ( n13990 , n13989 );
or ( n13991 , n13981 , n13990 );
not ( n13992 , n3764 );
and ( n13993 , n13992 , n4219 );
not ( n13994 , n4219 );
and ( n13995 , n13984 , n13985 );
xor ( n13996 , n13994 , n13995 );
and ( n13997 , n13996 , n3764 );
or ( n13998 , n13993 , n13997 );
not ( n13999 , n13998 );
not ( n14000 , n13999 );
or ( n14001 , n13991 , n14000 );
not ( n14002 , n3764 );
and ( n14003 , n14002 , n4209 );
not ( n14004 , n4209 );
and ( n14005 , n13994 , n13995 );
xor ( n14006 , n14004 , n14005 );
and ( n14007 , n14006 , n3764 );
or ( n14008 , n14003 , n14007 );
not ( n14009 , n14008 );
not ( n14010 , n14009 );
or ( n14011 , n14001 , n14010 );
not ( n14012 , n3764 );
and ( n14013 , n14012 , n4199 );
not ( n14014 , n4199 );
and ( n14015 , n14004 , n14005 );
xor ( n14016 , n14014 , n14015 );
and ( n14017 , n14016 , n3764 );
or ( n14018 , n14013 , n14017 );
not ( n14019 , n14018 );
not ( n14020 , n14019 );
or ( n14021 , n14011 , n14020 );
not ( n14022 , n3764 );
and ( n14023 , n14022 , n4189 );
not ( n14024 , n4189 );
and ( n14025 , n14014 , n14015 );
xor ( n14026 , n14024 , n14025 );
and ( n14027 , n14026 , n3764 );
or ( n14028 , n14023 , n14027 );
not ( n14029 , n14028 );
not ( n14030 , n14029 );
or ( n14031 , n14021 , n14030 );
not ( n14032 , n3764 );
and ( n14033 , n14032 , n4179 );
not ( n14034 , n4179 );
and ( n14035 , n14024 , n14025 );
xor ( n14036 , n14034 , n14035 );
and ( n14037 , n14036 , n3764 );
or ( n14038 , n14033 , n14037 );
not ( n14039 , n14038 );
not ( n14040 , n14039 );
or ( n14041 , n14031 , n14040 );
not ( n14042 , n3764 );
and ( n14043 , n14042 , n4169 );
not ( n14044 , n4169 );
and ( n14045 , n14034 , n14035 );
xor ( n14046 , n14044 , n14045 );
and ( n14047 , n14046 , n3764 );
or ( n14048 , n14043 , n14047 );
not ( n14049 , n14048 );
not ( n14050 , n14049 );
or ( n14051 , n14041 , n14050 );
not ( n14052 , n3764 );
and ( n14053 , n14052 , n4159 );
not ( n14054 , n4159 );
and ( n14055 , n14044 , n14045 );
xor ( n14056 , n14054 , n14055 );
and ( n14057 , n14056 , n3764 );
or ( n14058 , n14053 , n14057 );
not ( n14059 , n14058 );
not ( n14060 , n14059 );
or ( n14061 , n14051 , n14060 );
not ( n14062 , n3764 );
and ( n14063 , n14062 , n4149 );
not ( n14064 , n4149 );
and ( n14065 , n14054 , n14055 );
xor ( n14066 , n14064 , n14065 );
and ( n14067 , n14066 , n3764 );
or ( n14068 , n14063 , n14067 );
not ( n14069 , n14068 );
not ( n14070 , n14069 );
or ( n14071 , n14061 , n14070 );
not ( n14072 , n3764 );
and ( n14073 , n14072 , n4139 );
not ( n14074 , n4139 );
and ( n14075 , n14064 , n14065 );
xor ( n14076 , n14074 , n14075 );
and ( n14077 , n14076 , n3764 );
or ( n14078 , n14073 , n14077 );
not ( n14079 , n14078 );
not ( n14080 , n14079 );
or ( n14081 , n14071 , n14080 );
not ( n14082 , n3764 );
and ( n14083 , n14082 , n4129 );
not ( n14084 , n4129 );
and ( n14085 , n14074 , n14075 );
xor ( n14086 , n14084 , n14085 );
and ( n14087 , n14086 , n3764 );
or ( n14088 , n14083 , n14087 );
not ( n14089 , n14088 );
not ( n14090 , n14089 );
or ( n14091 , n14081 , n14090 );
not ( n14092 , n3764 );
and ( n14093 , n14092 , n4119 );
not ( n14094 , n4119 );
and ( n14095 , n14084 , n14085 );
xor ( n14096 , n14094 , n14095 );
and ( n14097 , n14096 , n3764 );
or ( n14098 , n14093 , n14097 );
not ( n14099 , n14098 );
not ( n14100 , n14099 );
or ( n14101 , n14091 , n14100 );
not ( n14102 , n3764 );
and ( n14103 , n14102 , n4109 );
not ( n14104 , n4109 );
and ( n14105 , n14094 , n14095 );
xor ( n14106 , n14104 , n14105 );
and ( n14107 , n14106 , n3764 );
or ( n14108 , n14103 , n14107 );
not ( n14109 , n14108 );
not ( n14110 , n14109 );
or ( n14111 , n14101 , n14110 );
not ( n14112 , n3764 );
and ( n14113 , n14112 , n4099 );
not ( n14114 , n4099 );
and ( n14115 , n14104 , n14105 );
xor ( n14116 , n14114 , n14115 );
and ( n14117 , n14116 , n3764 );
or ( n14118 , n14113 , n14117 );
not ( n14119 , n14118 );
not ( n14120 , n14119 );
or ( n14121 , n14111 , n14120 );
not ( n14122 , n3764 );
and ( n14123 , n14122 , n4089 );
not ( n14124 , n4089 );
and ( n14125 , n14114 , n14115 );
xor ( n14126 , n14124 , n14125 );
and ( n14127 , n14126 , n3764 );
or ( n14128 , n14123 , n14127 );
not ( n14129 , n14128 );
not ( n14130 , n14129 );
or ( n14131 , n14121 , n14130 );
not ( n14132 , n3764 );
and ( n14133 , n14132 , n4079 );
not ( n14134 , n4079 );
and ( n14135 , n14124 , n14125 );
xor ( n14136 , n14134 , n14135 );
and ( n14137 , n14136 , n3764 );
or ( n14138 , n14133 , n14137 );
not ( n14139 , n14138 );
not ( n14140 , n14139 );
or ( n14141 , n14131 , n14140 );
and ( n14142 , n14141 , n3764 );
not ( n14143 , n14142 );
and ( n14144 , n14143 , n13951 );
xor ( n14145 , n13951 , n3764 );
xor ( n14146 , n14145 , n3764 );
and ( n14147 , n14146 , n14142 );
or ( n14148 , n14144 , n14147 );
xor ( n14149 , n14148 , n13947 );
and ( n14150 , n14149 , n5287 );
or ( n14151 , n5154 , n5152 );
and ( n14152 , n5490 , n14151 );
or ( n14153 , n13949 , n14150 , n14152 );
not ( n14154 , n14153 );
not ( n14155 , n14154 );
buf ( n14156 , n14155 );
and ( n14157 , n14156 , n3259 );
or ( n14158 , n13746 , n14157 );
and ( n14159 , n13722 , n14158 );
and ( n14160 , n13743 , n3066 );
or ( n14161 , n14159 , n14160 );
and ( n14162 , n14161 , n2422 );
buf ( n14163 , n4245 );
not ( n14164 , n14163 );
not ( n14165 , n14164 );
buf ( n14166 , n14165 );
and ( n14167 , n14166 , n2428 );
or ( n14168 , n14162 , n14167 );
buf ( n14169 , n14168 );
buf ( n14170 , n2424 );
buf ( n14171 , n2281 );
buf ( n14172 , n2280 );
not ( n14173 , n3066 );
not ( n14174 , n3259 );
and ( n14175 , n2346 , n12991 );
not ( n14176 , n13313 );
and ( n14177 , n14176 , n13119 );
xor ( n14178 , n13119 , n13084 );
and ( n14179 , n13727 , n13728 );
xor ( n14180 , n14178 , n14179 );
and ( n14181 , n14180 , n13313 );
or ( n14182 , n14177 , n14181 );
and ( n14183 , n14182 , n5289 );
not ( n14184 , n13641 );
and ( n14185 , n14184 , n13447 );
xor ( n14186 , n13447 , n13412 );
and ( n14187 , n13735 , n13736 );
xor ( n14188 , n14186 , n14187 );
and ( n14189 , n14188 , n13641 );
or ( n14190 , n14185 , n14189 );
and ( n14191 , n14190 , n5287 );
and ( n14192 , n5735 , n5152 );
and ( n14193 , n2346 , n5154 );
or ( n14194 , n14183 , n14191 , n14192 , n14193 );
and ( n14195 , n14194 , n13662 );
or ( n14196 , n14175 , n14195 );
and ( n14197 , n14174 , n14196 );
and ( n14198 , n2424 , n3259 );
or ( n14199 , n14197 , n14198 );
and ( n14200 , n14173 , n14199 );
and ( n14201 , n14194 , n3066 );
or ( n14202 , n14200 , n14201 );
and ( n14203 , n14202 , n2422 );
buf ( n14204 , n3945 );
not ( n14205 , n14204 );
not ( n14206 , n14205 );
buf ( n14207 , n14206 );
and ( n14208 , n14207 , n2428 );
or ( n14209 , n14203 , n14208 );
buf ( n14210 , n14209 );
buf ( n14211 , n2424 );
buf ( n14212 , n2281 );
buf ( n14213 , n2280 );
not ( n14214 , n3066 );
not ( n14215 , n3259 );
and ( n14216 , n2344 , n12991 );
not ( n14217 , n13313 );
and ( n14218 , n14217 , n13131 );
xor ( n14219 , n13131 , n13084 );
and ( n14220 , n14178 , n14179 );
xor ( n14221 , n14219 , n14220 );
and ( n14222 , n14221 , n13313 );
or ( n14223 , n14218 , n14222 );
and ( n14224 , n14223 , n5289 );
not ( n14225 , n13641 );
and ( n14226 , n14225 , n13459 );
xor ( n14227 , n13459 , n13412 );
and ( n14228 , n14186 , n14187 );
xor ( n14229 , n14227 , n14228 );
and ( n14230 , n14229 , n13641 );
or ( n14231 , n14226 , n14230 );
and ( n14232 , n14231 , n5287 );
and ( n14233 , n5725 , n5152 );
and ( n14234 , n2344 , n5154 );
or ( n14235 , n14224 , n14232 , n14233 , n14234 );
and ( n14236 , n14235 , n13662 );
or ( n14237 , n14216 , n14236 );
and ( n14238 , n14215 , n14237 );
buf ( n14239 , n14156 );
and ( n14240 , n14239 , n3259 );
or ( n14241 , n14238 , n14240 );
and ( n14242 , n14214 , n14241 );
and ( n14243 , n14235 , n3066 );
or ( n14244 , n14242 , n14243 );
and ( n14245 , n14244 , n2422 );
buf ( n14246 , n3940 );
not ( n14247 , n14246 );
not ( n14248 , n14247 );
buf ( n14249 , n14248 );
and ( n14250 , n14249 , n2428 );
or ( n14251 , n14245 , n14250 );
buf ( n14252 , n14251 );
buf ( n14253 , n2424 );
buf ( n14254 , n2281 );
buf ( n14255 , n2280 );
not ( n14256 , n3066 );
not ( n14257 , n3259 );
and ( n14258 , n2342 , n12991 );
not ( n14259 , n13313 );
and ( n14260 , n14259 , n13143 );
xor ( n14261 , n13143 , n13084 );
and ( n14262 , n14219 , n14220 );
xor ( n14263 , n14261 , n14262 );
and ( n14264 , n14263 , n13313 );
or ( n14265 , n14260 , n14264 );
and ( n14266 , n14265 , n5289 );
not ( n14267 , n13641 );
and ( n14268 , n14267 , n13471 );
xor ( n14269 , n13471 , n13412 );
and ( n14270 , n14227 , n14228 );
xor ( n14271 , n14269 , n14270 );
and ( n14272 , n14271 , n13641 );
or ( n14273 , n14268 , n14272 );
and ( n14274 , n14273 , n5287 );
and ( n14275 , n5715 , n5152 );
and ( n14276 , n2342 , n5154 );
or ( n14277 , n14266 , n14274 , n14275 , n14276 );
and ( n14278 , n14277 , n13662 );
or ( n14279 , n14258 , n14278 );
and ( n14280 , n14257 , n14279 );
and ( n14281 , n2424 , n3259 );
or ( n14282 , n14280 , n14281 );
and ( n14283 , n14256 , n14282 );
and ( n14284 , n14277 , n3066 );
or ( n14285 , n14283 , n14284 );
and ( n14286 , n14285 , n2422 );
buf ( n14287 , n3935 );
not ( n14288 , n14287 );
not ( n14289 , n14288 );
buf ( n14290 , n14289 );
and ( n14291 , n14290 , n2428 );
or ( n14292 , n14286 , n14291 );
buf ( n14293 , n14292 );
buf ( n14294 , n2424 );
buf ( n14295 , n2281 );
buf ( n14296 , n2280 );
not ( n14297 , n3066 );
not ( n14298 , n3259 );
and ( n14299 , n2340 , n12991 );
not ( n14300 , n13313 );
and ( n14301 , n14300 , n13155 );
xor ( n14302 , n13155 , n13084 );
and ( n14303 , n14261 , n14262 );
xor ( n14304 , n14302 , n14303 );
and ( n14305 , n14304 , n13313 );
or ( n14306 , n14301 , n14305 );
and ( n14307 , n14306 , n5289 );
not ( n14308 , n13641 );
and ( n14309 , n14308 , n13483 );
or ( n14310 , n13483 , n13412 );
and ( n14311 , n14269 , n14270 );
xor ( n14312 , n14310 , n14311 );
and ( n14313 , n14312 , n13641 );
or ( n14314 , n14309 , n14313 );
and ( n14315 , n14314 , n5287 );
and ( n14316 , n5705 , n5152 );
and ( n14317 , n2340 , n5154 );
or ( n14318 , n14307 , n14315 , n14316 , n14317 );
and ( n14319 , n14318 , n13662 );
or ( n14320 , n14299 , n14319 );
and ( n14321 , n14298 , n14320 );
and ( n14322 , n2424 , n3259 );
or ( n14323 , n14321 , n14322 );
and ( n14324 , n14297 , n14323 );
and ( n14325 , n14318 , n3066 );
or ( n14326 , n14324 , n14325 );
and ( n14327 , n14326 , n2422 );
buf ( n14328 , n3930 );
not ( n14329 , n14328 );
not ( n14330 , n14329 );
buf ( n14331 , n14330 );
and ( n14332 , n14331 , n2428 );
or ( n14333 , n14327 , n14332 );
buf ( n14334 , n14333 );
buf ( n14335 , n2424 );
buf ( n14336 , n2281 );
buf ( n14337 , n2280 );
not ( n14338 , n3066 );
not ( n14339 , n3259 );
and ( n14340 , n2338 , n12991 );
not ( n14341 , n13313 );
and ( n14342 , n14341 , n13167 );
xor ( n14343 , n13167 , n13084 );
and ( n14344 , n14302 , n14303 );
xor ( n14345 , n14343 , n14344 );
and ( n14346 , n14345 , n13313 );
or ( n14347 , n14342 , n14346 );
and ( n14348 , n14347 , n5289 );
not ( n14349 , n13641 );
and ( n14350 , n14349 , n13495 );
xor ( n14351 , n13495 , n13412 );
and ( n14352 , n14310 , n14311 );
xor ( n14353 , n14351 , n14352 );
and ( n14354 , n14353 , n13641 );
or ( n14355 , n14350 , n14354 );
and ( n14356 , n14355 , n5287 );
and ( n14357 , n5695 , n5152 );
and ( n14358 , n2338 , n5154 );
or ( n14359 , n14348 , n14356 , n14357 , n14358 );
and ( n14360 , n14359 , n13662 );
or ( n14361 , n14340 , n14360 );
and ( n14362 , n14339 , n14361 );
and ( n14363 , n2424 , n3259 );
or ( n14364 , n14362 , n14363 );
and ( n14365 , n14338 , n14364 );
and ( n14366 , n14359 , n3066 );
or ( n14367 , n14365 , n14366 );
and ( n14368 , n14367 , n2422 );
buf ( n14369 , n3925 );
not ( n14370 , n14369 );
not ( n14371 , n14370 );
buf ( n14372 , n14371 );
and ( n14373 , n14372 , n2428 );
or ( n14374 , n14368 , n14373 );
buf ( n14375 , n14374 );
buf ( n14376 , n2424 );
buf ( n14377 , n2281 );
buf ( n14378 , n2280 );
not ( n14379 , n3066 );
not ( n14380 , n3259 );
and ( n14381 , n2336 , n12991 );
not ( n14382 , n13313 );
and ( n14383 , n14382 , n13179 );
xor ( n14384 , n13179 , n13084 );
and ( n14385 , n14343 , n14344 );
xor ( n14386 , n14384 , n14385 );
and ( n14387 , n14386 , n13313 );
or ( n14388 , n14383 , n14387 );
and ( n14389 , n14388 , n5289 );
not ( n14390 , n13641 );
and ( n14391 , n14390 , n13507 );
xor ( n14392 , n13507 , n13412 );
and ( n14393 , n14351 , n14352 );
xor ( n14394 , n14392 , n14393 );
and ( n14395 , n14394 , n13641 );
or ( n14396 , n14391 , n14395 );
and ( n14397 , n14396 , n5287 );
and ( n14398 , n5685 , n5152 );
and ( n14399 , n2336 , n5154 );
or ( n14400 , n14389 , n14397 , n14398 , n14399 );
and ( n14401 , n14400 , n13662 );
or ( n14402 , n14381 , n14401 );
and ( n14403 , n14380 , n14402 );
and ( n14404 , n2424 , n3259 );
or ( n14405 , n14403 , n14404 );
and ( n14406 , n14379 , n14405 );
and ( n14407 , n14400 , n3066 );
or ( n14408 , n14406 , n14407 );
and ( n14409 , n14408 , n2422 );
buf ( n14410 , n3920 );
not ( n14411 , n14410 );
not ( n14412 , n14411 );
buf ( n14413 , n14412 );
and ( n14414 , n14413 , n2428 );
or ( n14415 , n14409 , n14414 );
buf ( n14416 , n14415 );
buf ( n14417 , n2424 );
buf ( n14418 , n2281 );
buf ( n14419 , n2280 );
not ( n14420 , n3066 );
not ( n14421 , n3259 );
and ( n14422 , n2334 , n12991 );
not ( n14423 , n13313 );
and ( n14424 , n14423 , n13191 );
xor ( n14425 , n13191 , n13084 );
and ( n14426 , n14384 , n14385 );
xor ( n14427 , n14425 , n14426 );
and ( n14428 , n14427 , n13313 );
or ( n14429 , n14424 , n14428 );
and ( n14430 , n14429 , n5289 );
not ( n14431 , n13641 );
and ( n14432 , n14431 , n13519 );
xor ( n14433 , n13519 , n13412 );
and ( n14434 , n14392 , n14393 );
xor ( n14435 , n14433 , n14434 );
and ( n14436 , n14435 , n13641 );
or ( n14437 , n14432 , n14436 );
and ( n14438 , n14437 , n5287 );
and ( n14439 , n5675 , n5152 );
and ( n14440 , n2334 , n5154 );
or ( n14441 , n14430 , n14438 , n14439 , n14440 );
and ( n14442 , n14441 , n13662 );
or ( n14443 , n14422 , n14442 );
and ( n14444 , n14421 , n14443 );
and ( n14445 , n2424 , n3259 );
or ( n14446 , n14444 , n14445 );
and ( n14447 , n14420 , n14446 );
and ( n14448 , n14441 , n3066 );
or ( n14449 , n14447 , n14448 );
and ( n14450 , n14449 , n2422 );
buf ( n14451 , n3915 );
not ( n14452 , n14451 );
not ( n14453 , n14452 );
buf ( n14454 , n14453 );
and ( n14455 , n14454 , n2428 );
or ( n14456 , n14450 , n14455 );
buf ( n14457 , n14456 );
buf ( n14458 , n2424 );
buf ( n14459 , n2281 );
buf ( n14460 , n2280 );
not ( n14461 , n3066 );
not ( n14462 , n3259 );
and ( n14463 , n2332 , n12991 );
not ( n14464 , n13313 );
and ( n14465 , n14464 , n13203 );
xor ( n14466 , n13203 , n13084 );
and ( n14467 , n14425 , n14426 );
xor ( n14468 , n14466 , n14467 );
and ( n14469 , n14468 , n13313 );
or ( n14470 , n14465 , n14469 );
and ( n14471 , n14470 , n5289 );
not ( n14472 , n13641 );
and ( n14473 , n14472 , n13531 );
xor ( n14474 , n13531 , n13412 );
and ( n14475 , n14433 , n14434 );
or ( n14476 , n14474 , n14475 );
and ( n14477 , n14476 , n13641 );
or ( n14478 , n14473 , n14477 );
and ( n14479 , n14478 , n5287 );
and ( n14480 , n5665 , n5152 );
and ( n14481 , n2332 , n5154 );
or ( n14482 , n14471 , n14479 , n14480 , n14481 );
and ( n14483 , n14482 , n13662 );
or ( n14484 , n14463 , n14483 );
and ( n14485 , n14462 , n14484 );
and ( n14486 , n2424 , n3259 );
or ( n14487 , n14485 , n14486 );
and ( n14488 , n14461 , n14487 );
and ( n14489 , n14482 , n3066 );
or ( n14490 , n14488 , n14489 );
and ( n14491 , n14490 , n2422 );
buf ( n14492 , n3910 );
not ( n14493 , n14492 );
not ( n14494 , n14493 );
buf ( n14495 , n14494 );
and ( n14496 , n14495 , n2428 );
or ( n14497 , n14491 , n14496 );
buf ( n14498 , n14497 );
buf ( n14499 , n2424 );
buf ( n14500 , n2281 );
buf ( n14501 , n2280 );
not ( n14502 , n3066 );
not ( n14503 , n3259 );
and ( n14504 , n2330 , n12991 );
not ( n14505 , n13313 );
and ( n14506 , n14505 , n13215 );
xor ( n14507 , n13215 , n13084 );
and ( n14508 , n14466 , n14467 );
xor ( n14509 , n14507 , n14508 );
and ( n14510 , n14509 , n13313 );
or ( n14511 , n14506 , n14510 );
and ( n14512 , n14511 , n5289 );
not ( n14513 , n13641 );
and ( n14514 , n14513 , n13543 );
xor ( n14515 , n13543 , n13412 );
and ( n14516 , n14474 , n14475 );
xor ( n14517 , n14515 , n14516 );
and ( n14518 , n14517 , n13641 );
or ( n14519 , n14514 , n14518 );
and ( n14520 , n14519 , n5287 );
and ( n14521 , n5655 , n5152 );
and ( n14522 , n2330 , n5154 );
or ( n14523 , n14512 , n14520 , n14521 , n14522 );
and ( n14524 , n14523 , n13662 );
or ( n14525 , n14504 , n14524 );
and ( n14526 , n14503 , n14525 );
and ( n14527 , n2424 , n3259 );
or ( n14528 , n14526 , n14527 );
and ( n14529 , n14502 , n14528 );
and ( n14530 , n14523 , n3066 );
or ( n14531 , n14529 , n14530 );
and ( n14532 , n14531 , n2422 );
buf ( n14533 , n3905 );
not ( n14534 , n14533 );
not ( n14535 , n14534 );
buf ( n14536 , n14535 );
and ( n14537 , n14536 , n2428 );
or ( n14538 , n14532 , n14537 );
buf ( n14539 , n14538 );
buf ( n14540 , n2424 );
buf ( n14541 , n2281 );
buf ( n14542 , n2280 );
not ( n14543 , n3066 );
not ( n14544 , n3259 );
and ( n14545 , n2328 , n12991 );
not ( n14546 , n13313 );
and ( n14547 , n14546 , n13227 );
xor ( n14548 , n13227 , n13084 );
and ( n14549 , n14507 , n14508 );
xor ( n14550 , n14548 , n14549 );
and ( n14551 , n14550 , n13313 );
or ( n14552 , n14547 , n14551 );
and ( n14553 , n14552 , n5289 );
not ( n14554 , n13641 );
and ( n14555 , n14554 , n13555 );
xor ( n14556 , n13555 , n13412 );
and ( n14557 , n14515 , n14516 );
xor ( n14558 , n14556 , n14557 );
and ( n14559 , n14558 , n13641 );
or ( n14560 , n14555 , n14559 );
and ( n14561 , n14560 , n5287 );
and ( n14562 , n5645 , n5152 );
and ( n14563 , n2328 , n5154 );
or ( n14564 , n14553 , n14561 , n14562 , n14563 );
and ( n14565 , n14564 , n13662 );
or ( n14566 , n14545 , n14565 );
and ( n14567 , n14544 , n14566 );
and ( n14568 , n2424 , n3259 );
or ( n14569 , n14567 , n14568 );
and ( n14570 , n14543 , n14569 );
and ( n14571 , n14564 , n3066 );
or ( n14572 , n14570 , n14571 );
and ( n14573 , n14572 , n2422 );
buf ( n14574 , n3900 );
not ( n14575 , n14574 );
not ( n14576 , n14575 );
buf ( n14577 , n14576 );
and ( n14578 , n14577 , n2428 );
or ( n14579 , n14573 , n14578 );
buf ( n14580 , n14579 );
buf ( n14581 , n2424 );
buf ( n14582 , n2281 );
buf ( n14583 , n2280 );
not ( n14584 , n3066 );
not ( n14585 , n3259 );
and ( n14586 , n2326 , n12991 );
not ( n14587 , n13313 );
and ( n14588 , n14587 , n13239 );
xor ( n14589 , n13239 , n13084 );
and ( n14590 , n14548 , n14549 );
xor ( n14591 , n14589 , n14590 );
and ( n14592 , n14591 , n13313 );
or ( n14593 , n14588 , n14592 );
and ( n14594 , n14593 , n5289 );
not ( n14595 , n13641 );
and ( n14596 , n14595 , n13567 );
xor ( n14597 , n13567 , n13412 );
and ( n14598 , n14556 , n14557 );
xor ( n14599 , n14597 , n14598 );
and ( n14600 , n14599 , n13641 );
or ( n14601 , n14596 , n14600 );
and ( n14602 , n14601 , n5287 );
and ( n14603 , n5635 , n5152 );
and ( n14604 , n2326 , n5154 );
or ( n14605 , n14594 , n14602 , n14603 , n14604 );
and ( n14606 , n14605 , n13662 );
or ( n14607 , n14586 , n14606 );
and ( n14608 , n14585 , n14607 );
and ( n14609 , n2424 , n3259 );
or ( n14610 , n14608 , n14609 );
and ( n14611 , n14584 , n14610 );
and ( n14612 , n14605 , n3066 );
or ( n14613 , n14611 , n14612 );
and ( n14614 , n14613 , n2422 );
buf ( n14615 , n3895 );
not ( n14616 , n14615 );
not ( n14617 , n14616 );
buf ( n14618 , n14617 );
and ( n14619 , n14618 , n2428 );
or ( n14620 , n14614 , n14619 );
buf ( n14621 , n14620 );
buf ( n14622 , n2424 );
buf ( n14623 , n2281 );
buf ( n14624 , n2280 );
not ( n14625 , n3066 );
not ( n14626 , n3259 );
and ( n14627 , n2324 , n12991 );
not ( n14628 , n13313 );
and ( n14629 , n14628 , n13251 );
xor ( n14630 , n13251 , n13084 );
and ( n14631 , n14589 , n14590 );
xor ( n14632 , n14630 , n14631 );
and ( n14633 , n14632 , n13313 );
or ( n14634 , n14629 , n14633 );
and ( n14635 , n14634 , n5289 );
not ( n14636 , n13641 );
and ( n14637 , n14636 , n13579 );
xor ( n14638 , n13579 , n13412 );
and ( n14639 , n14597 , n14598 );
xor ( n14640 , n14638 , n14639 );
and ( n14641 , n14640 , n13641 );
or ( n14642 , n14637 , n14641 );
and ( n14643 , n14642 , n5287 );
and ( n14644 , n5625 , n5152 );
and ( n14645 , n2324 , n5154 );
or ( n14646 , n14635 , n14643 , n14644 , n14645 );
and ( n14647 , n14646 , n13662 );
or ( n14648 , n14627 , n14647 );
and ( n14649 , n14626 , n14648 );
and ( n14650 , n2424 , n3259 );
or ( n14651 , n14649 , n14650 );
and ( n14652 , n14625 , n14651 );
and ( n14653 , n14646 , n3066 );
or ( n14654 , n14652 , n14653 );
and ( n14655 , n14654 , n2422 );
buf ( n14656 , n3890 );
not ( n14657 , n14656 );
not ( n14658 , n14657 );
buf ( n14659 , n14658 );
and ( n14660 , n14659 , n2428 );
or ( n14661 , n14655 , n14660 );
buf ( n14662 , n14661 );
buf ( n14663 , n2424 );
buf ( n14664 , n2281 );
buf ( n14665 , n2280 );
not ( n14666 , n3066 );
not ( n14667 , n3259 );
and ( n14668 , n2322 , n12991 );
not ( n14669 , n13313 );
and ( n14670 , n14669 , n13263 );
xor ( n14671 , n13263 , n13084 );
and ( n14672 , n14630 , n14631 );
xor ( n14673 , n14671 , n14672 );
and ( n14674 , n14673 , n13313 );
or ( n14675 , n14670 , n14674 );
and ( n14676 , n14675 , n5289 );
not ( n14677 , n13641 );
and ( n14678 , n14677 , n13591 );
xor ( n14679 , n13591 , n13412 );
and ( n14680 , n14638 , n14639 );
xor ( n14681 , n14679 , n14680 );
and ( n14682 , n14681 , n13641 );
or ( n14683 , n14678 , n14682 );
and ( n14684 , n14683 , n5287 );
and ( n14685 , n5615 , n5152 );
and ( n14686 , n2322 , n5154 );
or ( n14687 , n14676 , n14684 , n14685 , n14686 );
and ( n14688 , n14687 , n13662 );
or ( n14689 , n14668 , n14688 );
and ( n14690 , n14667 , n14689 );
and ( n14691 , n2424 , n3259 );
or ( n14692 , n14690 , n14691 );
and ( n14693 , n14666 , n14692 );
and ( n14694 , n14687 , n3066 );
or ( n14695 , n14693 , n14694 );
and ( n14696 , n14695 , n2422 );
buf ( n14697 , n3885 );
not ( n14698 , n14697 );
not ( n14699 , n14698 );
buf ( n14700 , n14699 );
and ( n14701 , n14700 , n2428 );
or ( n14702 , n14696 , n14701 );
buf ( n14703 , n14702 );
buf ( n14704 , n2424 );
buf ( n14705 , n2281 );
buf ( n14706 , n2280 );
not ( n14707 , n3066 );
not ( n14708 , n3259 );
and ( n14709 , n2320 , n12991 );
not ( n14710 , n13313 );
and ( n14711 , n14710 , n13275 );
xor ( n14712 , n13275 , n13084 );
and ( n14713 , n14671 , n14672 );
xor ( n14714 , n14712 , n14713 );
and ( n14715 , n14714 , n13313 );
or ( n14716 , n14711 , n14715 );
and ( n14717 , n14716 , n5289 );
not ( n14718 , n13641 );
and ( n14719 , n14718 , n13603 );
xor ( n14720 , n13603 , n13412 );
and ( n14721 , n14679 , n14680 );
xor ( n14722 , n14720 , n14721 );
and ( n14723 , n14722 , n13641 );
or ( n14724 , n14719 , n14723 );
and ( n14725 , n14724 , n5287 );
and ( n14726 , n5605 , n5152 );
and ( n14727 , n2320 , n5154 );
or ( n14728 , n14717 , n14725 , n14726 , n14727 );
and ( n14729 , n14728 , n13662 );
or ( n14730 , n14709 , n14729 );
and ( n14731 , n14708 , n14730 );
and ( n14732 , n2424 , n3259 );
or ( n14733 , n14731 , n14732 );
and ( n14734 , n14707 , n14733 );
and ( n14735 , n14728 , n3066 );
or ( n14736 , n14734 , n14735 );
and ( n14737 , n14736 , n2422 );
buf ( n14738 , n3880 );
not ( n14739 , n14738 );
not ( n14740 , n14739 );
buf ( n14741 , n14740 );
and ( n14742 , n14741 , n2428 );
or ( n14743 , n14737 , n14742 );
buf ( n14744 , n14743 );
buf ( n14745 , n2424 );
buf ( n14746 , n2281 );
buf ( n14747 , n2280 );
not ( n14748 , n3066 );
not ( n14749 , n3259 );
and ( n14750 , n2318 , n12991 );
not ( n14751 , n13313 );
and ( n14752 , n14751 , n13287 );
xor ( n14753 , n13287 , n13084 );
and ( n14754 , n14712 , n14713 );
xor ( n14755 , n14753 , n14754 );
and ( n14756 , n14755 , n13313 );
or ( n14757 , n14752 , n14756 );
and ( n14758 , n14757 , n5289 );
not ( n14759 , n13641 );
and ( n14760 , n14759 , n13615 );
xor ( n14761 , n13615 , n13412 );
and ( n14762 , n14720 , n14721 );
xor ( n14763 , n14761 , n14762 );
and ( n14764 , n14763 , n13641 );
or ( n14765 , n14760 , n14764 );
and ( n14766 , n14765 , n5287 );
and ( n14767 , n5595 , n5152 );
and ( n14768 , n2318 , n5154 );
or ( n14769 , n14758 , n14766 , n14767 , n14768 );
and ( n14770 , n14769 , n13662 );
or ( n14771 , n14750 , n14770 );
and ( n14772 , n14749 , n14771 );
and ( n14773 , n2424 , n3259 );
or ( n14774 , n14772 , n14773 );
and ( n14775 , n14748 , n14774 );
and ( n14776 , n14769 , n3066 );
or ( n14777 , n14775 , n14776 );
and ( n14778 , n14777 , n2422 );
buf ( n14779 , n3875 );
not ( n14780 , n14779 );
not ( n14781 , n14780 );
buf ( n14782 , n14781 );
and ( n14783 , n14782 , n2428 );
or ( n14784 , n14778 , n14783 );
buf ( n14785 , n14784 );
buf ( n14786 , n2424 );
buf ( n14787 , n2281 );
buf ( n14788 , n2280 );
not ( n14789 , n3066 );
not ( n14790 , n3259 );
and ( n14791 , n2316 , n12991 );
not ( n14792 , n13313 );
and ( n14793 , n14792 , n13299 );
xor ( n14794 , n13299 , n13084 );
and ( n14795 , n14753 , n14754 );
xor ( n14796 , n14794 , n14795 );
and ( n14797 , n14796 , n13313 );
or ( n14798 , n14793 , n14797 );
and ( n14799 , n14798 , n5289 );
not ( n14800 , n13641 );
and ( n14801 , n14800 , n13627 );
xor ( n14802 , n13627 , n13412 );
and ( n14803 , n14761 , n14762 );
xor ( n14804 , n14802 , n14803 );
and ( n14805 , n14804 , n13641 );
or ( n14806 , n14801 , n14805 );
and ( n14807 , n14806 , n5287 );
and ( n14808 , n5585 , n5152 );
and ( n14809 , n2316 , n5154 );
or ( n14810 , n14799 , n14807 , n14808 , n14809 );
and ( n14811 , n14810 , n13662 );
or ( n14812 , n14791 , n14811 );
and ( n14813 , n14790 , n14812 );
and ( n14814 , n2424 , n3259 );
or ( n14815 , n14813 , n14814 );
and ( n14816 , n14789 , n14815 );
and ( n14817 , n14810 , n3066 );
or ( n14818 , n14816 , n14817 );
and ( n14819 , n14818 , n2422 );
buf ( n14820 , n3870 );
not ( n14821 , n14820 );
not ( n14822 , n14821 );
buf ( n14823 , n14822 );
and ( n14824 , n14823 , n2428 );
or ( n14825 , n14819 , n14824 );
buf ( n14826 , n14825 );
buf ( n14827 , n2424 );
buf ( n14828 , n2281 );
buf ( n14829 , n2280 );
not ( n14830 , n3066 );
not ( n14831 , n3259 );
and ( n14832 , n2314 , n12991 );
not ( n14833 , n13313 );
and ( n14834 , n14833 , n13311 );
xor ( n14835 , n13311 , n13084 );
and ( n14836 , n14794 , n14795 );
xor ( n14837 , n14835 , n14836 );
and ( n14838 , n14837 , n13313 );
or ( n14839 , n14834 , n14838 );
and ( n14840 , n14839 , n5289 );
not ( n14841 , n13641 );
and ( n14842 , n14841 , n13639 );
xor ( n14843 , n13639 , n13412 );
and ( n14844 , n14802 , n14803 );
xor ( n14845 , n14843 , n14844 );
and ( n14846 , n14845 , n13641 );
or ( n14847 , n14842 , n14846 );
and ( n14848 , n14847 , n5287 );
and ( n14849 , n5575 , n5152 );
and ( n14850 , n2314 , n5154 );
or ( n14851 , n14840 , n14848 , n14849 , n14850 );
and ( n14852 , n14851 , n13662 );
or ( n14853 , n14832 , n14852 );
and ( n14854 , n14831 , n14853 );
and ( n14855 , n2424 , n3259 );
or ( n14856 , n14854 , n14855 );
and ( n14857 , n14830 , n14856 );
and ( n14858 , n14851 , n3066 );
or ( n14859 , n14857 , n14858 );
and ( n14860 , n14859 , n2422 );
buf ( n14861 , n3865 );
not ( n14862 , n14861 );
not ( n14863 , n14862 );
buf ( n14864 , n14863 );
and ( n14865 , n14864 , n2428 );
or ( n14866 , n14860 , n14865 );
buf ( n14867 , n14866 );
buf ( n14868 , n2424 );
buf ( n14869 , n2281 );
buf ( n14870 , n2280 );
not ( n14871 , n3259 );
or ( n14872 , n3066 , n14871 );
not ( n14873 , n14872 );
and ( n14874 , n14873 , n3795 );
and ( n14875 , n2416 , n14872 );
or ( n14876 , n14874 , n14875 );
and ( n14877 , n14876 , n2422 );
and ( n14878 , n2416 , n2428 );
or ( n14879 , n14877 , n14878 );
buf ( n14880 , n14879 );
buf ( n14881 , n2424 );
buf ( n14882 , n2281 );
buf ( n14883 , n2280 );
not ( n14884 , n14872 );
and ( n14885 , n14884 , n3785 );
and ( n14886 , n2414 , n14872 );
or ( n14887 , n14885 , n14886 );
and ( n14888 , n14887 , n2422 );
and ( n14889 , n2414 , n2428 );
or ( n14890 , n14888 , n14889 );
buf ( n14891 , n14890 );
buf ( n14892 , n2424 );
buf ( n14893 , n2281 );
buf ( n14894 , n2280 );
not ( n14895 , n14872 );
and ( n14896 , n14895 , n4257 );
and ( n14897 , n2412 , n14872 );
or ( n14898 , n14896 , n14897 );
and ( n14899 , n14898 , n2422 );
and ( n14900 , n2412 , n2428 );
or ( n14901 , n14899 , n14900 );
buf ( n14902 , n14901 );
buf ( n14903 , n2424 );
buf ( n14904 , n2281 );
buf ( n14905 , n2280 );
not ( n14906 , n14872 );
and ( n14907 , n14906 , n4243 );
and ( n14908 , n2410 , n14872 );
or ( n14909 , n14907 , n14908 );
and ( n14910 , n14909 , n2422 );
and ( n14911 , n2410 , n2428 );
or ( n14912 , n14910 , n14911 );
buf ( n14913 , n14912 );
buf ( n14914 , n2424 );
buf ( n14915 , n2281 );
buf ( n14916 , n2280 );
not ( n14917 , n14872 );
and ( n14918 , n14917 , n4233 );
and ( n14919 , n2408 , n14872 );
or ( n14920 , n14918 , n14919 );
and ( n14921 , n14920 , n2422 );
and ( n14922 , n2408 , n2428 );
or ( n14923 , n14921 , n14922 );
buf ( n14924 , n14923 );
buf ( n14925 , n2424 );
buf ( n14926 , n2281 );
buf ( n14927 , n2280 );
not ( n14928 , n14872 );
and ( n14929 , n14928 , n4223 );
and ( n14930 , n2406 , n14872 );
or ( n14931 , n14929 , n14930 );
and ( n14932 , n14931 , n2422 );
and ( n14933 , n2406 , n2428 );
or ( n14934 , n14932 , n14933 );
buf ( n14935 , n14934 );
buf ( n14936 , n2424 );
buf ( n14937 , n2281 );
buf ( n14938 , n2280 );
not ( n14939 , n14872 );
and ( n14940 , n14939 , n4213 );
and ( n14941 , n2404 , n14872 );
or ( n14942 , n14940 , n14941 );
and ( n14943 , n14942 , n2422 );
and ( n14944 , n2404 , n2428 );
or ( n14945 , n14943 , n14944 );
buf ( n14946 , n14945 );
buf ( n14947 , n2424 );
buf ( n14948 , n2281 );
buf ( n14949 , n2280 );
not ( n14950 , n14872 );
and ( n14951 , n14950 , n4203 );
and ( n14952 , n2402 , n14872 );
or ( n14953 , n14951 , n14952 );
and ( n14954 , n14953 , n2422 );
and ( n14955 , n2402 , n2428 );
or ( n14956 , n14954 , n14955 );
buf ( n14957 , n14956 );
buf ( n14958 , n2424 );
buf ( n14959 , n2281 );
buf ( n14960 , n2280 );
not ( n14961 , n14872 );
and ( n14962 , n14961 , n4193 );
and ( n14963 , n2400 , n14872 );
or ( n14964 , n14962 , n14963 );
and ( n14965 , n14964 , n2422 );
and ( n14966 , n2400 , n2428 );
or ( n14967 , n14965 , n14966 );
buf ( n14968 , n14967 );
buf ( n14969 , n2424 );
buf ( n14970 , n2281 );
buf ( n14971 , n2280 );
not ( n14972 , n14872 );
and ( n14973 , n14972 , n4183 );
and ( n14974 , n2398 , n14872 );
or ( n14975 , n14973 , n14974 );
and ( n14976 , n14975 , n2422 );
and ( n14977 , n2398 , n2428 );
or ( n14978 , n14976 , n14977 );
buf ( n14979 , n14978 );
buf ( n14980 , n2424 );
buf ( n14981 , n2281 );
buf ( n14982 , n2280 );
not ( n14983 , n14872 );
and ( n14984 , n14983 , n4173 );
and ( n14985 , n2396 , n14872 );
or ( n14986 , n14984 , n14985 );
and ( n14987 , n14986 , n2422 );
and ( n14988 , n2396 , n2428 );
or ( n14989 , n14987 , n14988 );
buf ( n14990 , n14989 );
buf ( n14991 , n2424 );
buf ( n14992 , n2281 );
buf ( n14993 , n2280 );
not ( n14994 , n14872 );
and ( n14995 , n14994 , n4163 );
and ( n14996 , n2394 , n14872 );
or ( n14997 , n14995 , n14996 );
and ( n14998 , n14997 , n2422 );
and ( n14999 , n2394 , n2428 );
or ( n15000 , n14998 , n14999 );
buf ( n15001 , n15000 );
buf ( n15002 , n2424 );
buf ( n15003 , n2281 );
buf ( n15004 , n2280 );
not ( n15005 , n14872 );
and ( n15006 , n15005 , n4153 );
and ( n15007 , n2392 , n14872 );
or ( n15008 , n15006 , n15007 );
and ( n15009 , n15008 , n2422 );
and ( n15010 , n2392 , n2428 );
or ( n15011 , n15009 , n15010 );
buf ( n15012 , n15011 );
buf ( n15013 , n2424 );
buf ( n15014 , n2281 );
buf ( n15015 , n2280 );
not ( n15016 , n14872 );
and ( n15017 , n15016 , n4143 );
and ( n15018 , n2390 , n14872 );
or ( n15019 , n15017 , n15018 );
and ( n15020 , n15019 , n2422 );
and ( n15021 , n2390 , n2428 );
or ( n15022 , n15020 , n15021 );
buf ( n15023 , n15022 );
buf ( n15024 , n2424 );
buf ( n15025 , n2281 );
buf ( n15026 , n2280 );
not ( n15027 , n14872 );
and ( n15028 , n15027 , n4133 );
and ( n15029 , n2388 , n14872 );
or ( n15030 , n15028 , n15029 );
and ( n15031 , n15030 , n2422 );
and ( n15032 , n2388 , n2428 );
or ( n15033 , n15031 , n15032 );
buf ( n15034 , n15033 );
buf ( n15035 , n2424 );
buf ( n15036 , n2281 );
buf ( n15037 , n2280 );
not ( n15038 , n14872 );
and ( n15039 , n15038 , n4123 );
and ( n15040 , n2386 , n14872 );
or ( n15041 , n15039 , n15040 );
and ( n15042 , n15041 , n2422 );
and ( n15043 , n2386 , n2428 );
or ( n15044 , n15042 , n15043 );
buf ( n15045 , n15044 );
buf ( n15046 , n2424 );
buf ( n15047 , n2281 );
buf ( n15048 , n2280 );
not ( n15049 , n14872 );
and ( n15050 , n15049 , n4113 );
and ( n15051 , n2384 , n14872 );
or ( n15052 , n15050 , n15051 );
and ( n15053 , n15052 , n2422 );
and ( n15054 , n2384 , n2428 );
or ( n15055 , n15053 , n15054 );
buf ( n15056 , n15055 );
buf ( n15057 , n2424 );
buf ( n15058 , n2281 );
buf ( n15059 , n2280 );
not ( n15060 , n14872 );
and ( n15061 , n15060 , n4103 );
and ( n15062 , n2382 , n14872 );
or ( n15063 , n15061 , n15062 );
and ( n15064 , n15063 , n2422 );
and ( n15065 , n2382 , n2428 );
or ( n15066 , n15064 , n15065 );
buf ( n15067 , n15066 );
buf ( n15068 , n2424 );
buf ( n15069 , n2281 );
buf ( n15070 , n2280 );
not ( n15071 , n14872 );
and ( n15072 , n15071 , n4093 );
and ( n15073 , n2380 , n14872 );
or ( n15074 , n15072 , n15073 );
and ( n15075 , n15074 , n2422 );
and ( n15076 , n2380 , n2428 );
or ( n15077 , n15075 , n15076 );
buf ( n15078 , n15077 );
buf ( n15079 , n2424 );
buf ( n15080 , n2281 );
buf ( n15081 , n2280 );
not ( n15082 , n14872 );
and ( n15083 , n15082 , n4083 );
and ( n15084 , n2378 , n14872 );
or ( n15085 , n15083 , n15084 );
and ( n15086 , n15085 , n2422 );
and ( n15087 , n2378 , n2428 );
or ( n15088 , n15086 , n15087 );
buf ( n15089 , n15088 );
buf ( n15090 , n2424 );
buf ( n15091 , n2281 );
buf ( n15092 , n2280 );
not ( n15093 , n14872 );
and ( n15094 , n15093 , n4073 );
and ( n15095 , n2376 , n14872 );
or ( n15096 , n15094 , n15095 );
and ( n15097 , n15096 , n2422 );
and ( n15098 , n2376 , n2428 );
or ( n15099 , n15097 , n15098 );
buf ( n15100 , n15099 );
buf ( n15101 , n2424 );
buf ( n15102 , n2281 );
buf ( n15103 , n2280 );
not ( n15104 , n14872 );
and ( n15105 , n15104 , n4063 );
and ( n15106 , n2374 , n14872 );
or ( n15107 , n15105 , n15106 );
and ( n15108 , n15107 , n2422 );
and ( n15109 , n2374 , n2428 );
or ( n15110 , n15108 , n15109 );
buf ( n15111 , n15110 );
buf ( n15112 , n2424 );
buf ( n15113 , n2281 );
buf ( n15114 , n2280 );
not ( n15115 , n14872 );
and ( n15116 , n15115 , n4053 );
and ( n15117 , n2372 , n14872 );
or ( n15118 , n15116 , n15117 );
and ( n15119 , n15118 , n2422 );
and ( n15120 , n2372 , n2428 );
or ( n15121 , n15119 , n15120 );
buf ( n15122 , n15121 );
buf ( n15123 , n2424 );
buf ( n15124 , n2281 );
buf ( n15125 , n2280 );
not ( n15126 , n14872 );
and ( n15127 , n15126 , n4043 );
and ( n15128 , n2370 , n14872 );
or ( n15129 , n15127 , n15128 );
and ( n15130 , n15129 , n2422 );
and ( n15131 , n2370 , n2428 );
or ( n15132 , n15130 , n15131 );
buf ( n15133 , n15132 );
buf ( n15134 , n2424 );
buf ( n15135 , n2281 );
buf ( n15136 , n2280 );
not ( n15137 , n14872 );
and ( n15138 , n15137 , n4033 );
and ( n15139 , n2368 , n14872 );
or ( n15140 , n15138 , n15139 );
and ( n15141 , n15140 , n2422 );
and ( n15142 , n2368 , n2428 );
or ( n15143 , n15141 , n15142 );
buf ( n15144 , n15143 );
buf ( n15145 , n2424 );
buf ( n15146 , n2281 );
buf ( n15147 , n2280 );
not ( n15148 , n14872 );
and ( n15149 , n15148 , n4023 );
and ( n15150 , n2366 , n14872 );
or ( n15151 , n15149 , n15150 );
and ( n15152 , n15151 , n2422 );
and ( n15153 , n2366 , n2428 );
or ( n15154 , n15152 , n15153 );
buf ( n15155 , n15154 );
buf ( n15156 , n2424 );
buf ( n15157 , n2281 );
buf ( n15158 , n2280 );
not ( n15159 , n14872 );
and ( n15160 , n15159 , n4013 );
and ( n15161 , n2364 , n14872 );
or ( n15162 , n15160 , n15161 );
and ( n15163 , n15162 , n2422 );
and ( n15164 , n2364 , n2428 );
or ( n15165 , n15163 , n15164 );
buf ( n15166 , n15165 );
buf ( n15167 , n2424 );
buf ( n15168 , n2281 );
buf ( n15169 , n2280 );
not ( n15170 , n14872 );
and ( n15171 , n15170 , n4003 );
and ( n15172 , n2362 , n14872 );
or ( n15173 , n15171 , n15172 );
and ( n15174 , n15173 , n2422 );
and ( n15175 , n2362 , n2428 );
or ( n15176 , n15174 , n15175 );
buf ( n15177 , n15176 );
buf ( n15178 , n2424 );
buf ( n15179 , n2281 );
buf ( n15180 , n2280 );
not ( n15181 , n14872 );
and ( n15182 , n15181 , n3993 );
and ( n15183 , n2360 , n14872 );
or ( n15184 , n15182 , n15183 );
and ( n15185 , n15184 , n2422 );
and ( n15186 , n2360 , n2428 );
or ( n15187 , n15185 , n15186 );
buf ( n15188 , n15187 );
buf ( n15189 , n2424 );
buf ( n15190 , n2281 );
buf ( n15191 , n2280 );
not ( n15192 , n14872 );
and ( n15193 , n15192 , n3983 );
and ( n15194 , n2358 , n14872 );
or ( n15195 , n15193 , n15194 );
and ( n15196 , n15195 , n2422 );
and ( n15197 , n2358 , n2428 );
or ( n15198 , n15196 , n15197 );
buf ( n15199 , n15198 );
buf ( n15200 , n2424 );
buf ( n15201 , n2281 );
buf ( n15202 , n2280 );
not ( n15203 , n14872 );
and ( n15204 , n15203 , n3819 );
and ( n15205 , n2356 , n14872 );
or ( n15206 , n15204 , n15205 );
and ( n15207 , n15206 , n2422 );
and ( n15208 , n2356 , n2428 );
or ( n15209 , n15207 , n15208 );
buf ( n15210 , n15209 );
buf ( n15211 , n2424 );
buf ( n15212 , n2281 );
buf ( n15213 , n2280 );
not ( n15214 , n14872 );
and ( n15215 , n15214 , n3770 );
and ( n15216 , n2354 , n14872 );
or ( n15217 , n15215 , n15216 );
and ( n15218 , n15217 , n2422 );
and ( n15219 , n2354 , n2428 );
or ( n15220 , n15218 , n15219 );
buf ( n15221 , n15220 );
buf ( n15222 , n2424 );
buf ( n15223 , n2281 );
buf ( n15224 , n2280 );
not ( n15225 , n3066 );
and ( n15226 , n5290 , n13662 );
not ( n15227 , n3259 );
and ( n15228 , n15226 , n15227 );
and ( n15229 , n15225 , n15228 );
and ( n15230 , n5290 , n3066 );
or ( n15231 , n15229 , n15230 );
and ( n15232 , n15231 , n2422 );
or ( n15233 , n15232 , n2428 );
buf ( n15234 , n15233 );
buf ( n15235 , n2424 );
buf ( n15236 , n2281 );
buf ( n15237 , n2280 );
not ( n15238 , n14872 );
and ( n15239 , n3259 , n15238 );
and ( n15240 , n15239 , n2422 );
buf ( n15241 , n15240 );
endmodule
