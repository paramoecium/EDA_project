module top ( PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D );
input PI_clock , PI_reset , n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , DFF_state_reg_Q , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , DFF_B_reg_Q , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , DFF_rd_reg_Q , DFF_wr_reg_Q;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , PO_rd , PO_wr , DFF_state_reg_S , DFF_state_reg_R , DFF_state_reg_CK , DFF_state_reg_D , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , DFF_B_reg_S , DFF_B_reg_R , DFF_B_reg_CK , DFF_B_reg_D , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , DFF_rd_reg_S , DFF_rd_reg_R , DFF_rd_reg_CK , DFF_rd_reg_D , DFF_wr_reg_S , DFF_wr_reg_R , DFF_wr_reg_CK , DFF_wr_reg_D;
wire n68634 , n68635 , n68636 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n68644 , n68645 , n68646 , n2508 , n2509 , n68649 , n68650 , n68651 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n68659 , n68660 , n68661 , n2523 , n2524 , n68664 , n68665 , n68666 , n2528 , n2529 , n68669 , n68670 , n2532 , n2533 , n2534 , n68674 , n68675 , n68676 , n2538 , n2539 , n68679 , n68680 , n68681 , n2543 , n2544 , n68684 , n68685 , n2547 , n2548 , n2549 , n68689 , n68690 , n68691 , n2553 , n2554 , n68694 , n68695 , n68696 , n2558 , n2559 , n68699 , n68700 , n2562 , n2563 , n2564 , n68704 , n68705 , n68706 , n2568 , n2569 , n68709 , n68710 , n68711 , n2573 , n2574 , n68714 , n68715 , n2577 , n2578 , n2579 , n68719 , n68720 , n68721 , n2583 , n2584 , n68724 , n68725 , n68726 , n2588 , n2589 , n68729 , n68730 , n2592 , n2593 , n2594 , n68734 , n68735 , n68736 , n2598 , n2599 , n68739 , n68740 , n68741 , n2603 , n2604 , n2605 , n2606 , n68746 , n68747 , n2609 , n68749 , n68750 , n68751 , n2613 , n68753 , n68754 , n68755 , n68756 , n2618 , n68758 , n68759 , n2621 , n2622 , n2623 , n2624 , n68764 , n68765 , n68766 , n2628 , n2629 , n68769 , n68770 , n68771 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n68779 , n68780 , n68781 , n2643 , n2644 , n68784 , n68785 , n68786 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n68794 , n68795 , n68796 , n2658 , n2659 , n68799 , n68800 , n68801 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n68809 , n68810 , n68811 , n2673 , n2674 , n68814 , n68815 , n68816 , n68817 , n68818 , n2680 , n2681 , n2682 , n68822 , n68823 , n68824 , n68825 , n68826 , n2688 , n2689 , n68829 , n68830 , n68831 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n68838 , n68839 , n68840 , n68841 , n2703 , n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n2710 , n68850 , n68851 , n68852 , n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 , n68863 , n68864 , n68865 , n68866 , n2728 , n68868 , n68869 , n68870 , n68871 , n68872 , n2734 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 , n2744 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n2753 , n68893 , n68894 , n68895 , n68896 , n2758 , n68898 , n68899 , n68900 , n68901 , n68902 , n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 , n2774 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 , n2784 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 , n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 , n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 , n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 , n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 , n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 , n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 , n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 , n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 , n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 , n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 , n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 , n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 , n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 , n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 , n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 , n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 , n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 , n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 , n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 , n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n3000 , n69140 , n69141 , n69142 , n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 , n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 , n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 , n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 , n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 , n69193 , n69194 , n69195 , n69196 , n3058 , n3059 , n69199 , n69200 , n69201 , n69202 , n69203 , n69204 , n3066 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 , n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 , n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 , n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 , n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 , n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 , n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 , n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 , n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 , n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 , n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 , n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 , n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 , n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 , n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 , n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 , n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 , n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 , n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 , n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 , n69413 , n69414 , n3276 , n69416 , n69417 , n69418 , n69419 , n69420 , n3282 , n69422 , n69423 , n69424 , n69425 , n69426 , n3288 , n69428 , n69429 , n69430 , n3292 , n69432 , n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n3301 , n69441 , n69442 , n3304 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 , n69453 , n69454 , n3316 , n69456 , n69457 , n69458 , n3320 , n69460 , n69461 , n69462 , n3324 , n69464 , n69465 , n3327 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 , n69473 , n69474 , n3336 , n69476 , n69477 , n69478 , n69479 , n69480 , n3342 , n69482 , n3344 , n69484 , n3346 , n69486 , n69487 , n69488 , n3350 , n69490 , n69491 , n69492 , n69493 , n69494 , n3356 , n69496 , n69497 , n3359 , n69499 , n69500 , n69501 , n69502 , n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 , n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 , n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 , n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 , n69543 , n3405 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n3412 , n69552 , n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 , n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 , n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n3442 , n69582 , n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n3450 , n69590 , n69591 , n69592 , n3454 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 , n69603 , n69604 , n3466 , n69606 , n69607 , n69608 , n3470 , n69610 , n69611 , n69612 , n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n69627 , n3489 , n69629 , n69630 , n69631 , n69632 , n69633 , n69634 , n69635 , n69636 , n3498 , n69638 , n69639 , n69640 , n69641 , n69642 , n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n3510 , n69650 , n69651 , n69652 , n3514 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 , n69663 , n69664 , n69665 , n69666 , n69667 , n3529 , n69669 , n69670 , n69671 , n69672 , n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 , n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n3552 , n69692 , n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n3561 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n3569 , n69709 , n69710 , n69711 , n69712 , n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n3580 , n69720 , n69721 , n69722 , n3584 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n3591 , n69731 , n69732 , n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 , n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 , n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n3620 , n69760 , n69761 , n69762 , n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 , n69773 , n69774 , n3636 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 , n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 , n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 , n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 , n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 , n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 , n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 , n69843 , n69844 , n69845 , n3707 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 , n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n3721 , n69861 , n69862 , n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 , n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 , n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 , n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n3771 , n69911 , n69912 , n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 , n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 , n69933 , n69934 , n69935 , n69936 , n69937 , n3799 , n69939 , n69940 , n69941 , n69942 , n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 , n69953 , n3815 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 , n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 , n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 , n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 , n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 , n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 , n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 , n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 , n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 , n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 , n70053 , n3915 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 , n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 , n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 , n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 , n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 , n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 , n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 , n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 , n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 , n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 , n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 , n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 , n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 , n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 , n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 , n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 , n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 , n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 , n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 , n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 , n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 , n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 , n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 , n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 , n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 , n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 , n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 , n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 , n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 , n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 , n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 , n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 , n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 , n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 , n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 , n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 , n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 , n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 , n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 , n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 , n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 , n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 , n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 , n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 , n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n4769 , n4770 , n70910 , n70911 , n70912 , n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 , n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 , n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 , n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 , n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 , n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 , n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 , n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 , n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 , n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 , n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n4881 , n71021 , n71022 , n4884 , n4885 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 , n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 , n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 , n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 , n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 , n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 , n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 , n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 , n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 , n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 , n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 , n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 , n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 , n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 , n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n5071 , n5072 , n71212 , n5074 , n5075 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 , n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 , n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 , n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 , n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 , n71263 , n71264 , n71265 , n71266 , n5128 , n71268 , n71269 , n71270 , n5132 , n71272 , n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 , n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 , n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 , n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 , n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 , n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 , n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 , n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 , n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 , n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 , n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 , n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 , n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 , n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n5300 , n71440 , n71441 , n71442 , n5304 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 , n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 , n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 , n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 , n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 , n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 , n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 , n5374 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 , n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 , n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 , n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 , n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 , n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 , n71573 , n71574 , n71575 , n71576 , n71577 , n5439 , n5440 , n71580 , n71581 , n71582 , n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 , n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 , n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 , n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 , n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 , n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 , n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 , n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 , n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 , n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 , n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 , n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 , n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 , n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n5582 , n71722 , n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n5591 , n5592 , n71732 , n5594 , n5595 , n71735 , n71736 , n71737 , n71738 , n71739 , n5601 , n71741 , n71742 , n5604 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 , n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 , n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n5631 , n71771 , n71772 , n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 , n5644 , n5645 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 , n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 , n5664 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 , n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n5681 , n5682 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 , n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n5701 , n5702 , n71842 , n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 , n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 , n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 , n5734 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n5742 , n71882 , n71883 , n5745 , n71885 , n71886 , n71887 , n71888 , n71889 , n5751 , n5752 , n71892 , n5754 , n5755 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 , n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 , n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 , n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 , n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 , n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 , n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 , n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 , n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 , n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 , n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 , n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 , n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 , n72023 , n72024 , n72025 , n72026 , n72027 , n5889 , n72029 , n72030 , n72031 , n72032 , n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 , n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 , n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 , n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 , n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 , n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 , n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 , n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 , n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 , n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 , n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 , n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 , n72153 , n72154 , n72155 , n6017 , n72157 , n72158 , n72159 , n6021 , n72161 , n72162 , n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 , n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 , n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 , n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 , n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n6077 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 , n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 , n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 , n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 , n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 , n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 , n72273 , n72274 , n6136 , n6137 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 , n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 , n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 , n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 , n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 , n6184 , n6185 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 , n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 , n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 , n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 , n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 , n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 , n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 , n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 , n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 , n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 , n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 , n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 , n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 , n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 , n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 , n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 , n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 , n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 , n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 , n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 , n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 , n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 , n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 , n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 , n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 , n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 , n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 , n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 , n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 , n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 , n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 , n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 , n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 , n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 , n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 , n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 , n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 , n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 , n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 , n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 , n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 , n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 , n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 , n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 , n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 , n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 , n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 , n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 , n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 , n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 , n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 , n72833 , n72834 , n6696 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 , n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 , n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 , n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 , n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 , n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 , n72913 , n72914 , n6776 , n6777 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 , n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 , n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 , n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 , n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 , n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 , n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 , n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n6852 , n72992 , n72993 , n72994 , n6856 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 , n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 , n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 , n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 , n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 , n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 , n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 , n73063 , n73064 , n6926 , n6927 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 , n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 , n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 , n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 , n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 , n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 , n73123 , n73124 , n73125 , n6987 , n73127 , n73128 , n73129 , n6991 , n73131 , n73132 , n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 , n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 , n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 , n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 , n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 , n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 , n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 , n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 , n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 , n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 , n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 , n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 , n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 , n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 , n73273 , n73274 , n73275 , n73276 , n73277 , n7139 , n73279 , n73280 , n73281 , n73282 , n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 , n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 , n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 , n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 , n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 , n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n7207 , n7208 , n73348 , n73349 , n73350 , n73351 , n73352 , n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 , n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 , n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 , n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 , n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 , n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 , n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 , n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 , n73443 , n7305 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 , n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 , n73463 , n73464 , n73465 , n7327 , n7328 , n73468 , n73469 , n73470 , n73471 , n73472 , n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 , n73483 , n73484 , n73485 , n73486 , n73487 , n7349 , n7350 , n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n73526 , n7388 , n7389 , n73529 , n7391 , n7392 , n73532 , n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 , n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 , n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 , n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 , n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 , n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 , n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 , n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 , n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 , n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 , n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 , n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 , n73673 , n73674 , n7536 , n7537 , n73677 , n7539 , n7540 , n73680 , n73681 , n73682 , n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 , n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 , n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 , n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 , n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 , n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 , n73753 , n73754 , n73755 , n73756 , n73757 , n7619 , n73759 , n73760 , n7622 , n7623 , n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 , n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n7640 , n7641 , n73781 , n73782 , n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 , n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 , n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 , n73813 , n73814 , n7676 , n7677 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 , n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n7692 , n7693 , n73833 , n73834 , n7696 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 , n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 , n7714 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 , n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 , n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 , n73883 , n73884 , n73885 , n73886 , n73887 , n7749 , n7750 , n73890 , n73891 , n73892 , n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 , n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 , n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 , n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n7793 , n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 , n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 , n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 , n73963 , n73964 , n73965 , n73966 , n73967 , n7829 , n7830 , n73970 , n7832 , n7833 , n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 , n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 , n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 , n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 , n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n7920 , n7921 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 , n74073 , n74074 , n7936 , n7937 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 , n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n7953 , n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 , n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n7971 , n7972 , n74112 , n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 , n74123 , n74124 , n74125 , n74126 , n7988 , n7989 , n74129 , n74130 , n7992 , n74132 , n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 , n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n8010 , n8011 , n74151 , n74152 , n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 , n74163 , n74164 , n8026 , n8027 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 , n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 , n74183 , n8045 , n8046 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 , n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 , n74203 , n74204 , n74205 , n8067 , n8068 , n74208 , n74209 , n74210 , n74211 , n74212 , n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 , n8084 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 , n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 , n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 , n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 , n74263 , n74264 , n8126 , n8127 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 , n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n8142 , n8143 , n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 , n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n8163 , n8164 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 , n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 , n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 , n74333 , n74334 , n74335 , n74336 , n74337 , n8199 , n74339 , n8201 , n8202 , n74342 , n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 , n74353 , n74354 , n74355 , n8217 , n74357 , n74358 , n74359 , n8221 , n74361 , n74362 , n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 , n74373 , n74374 , n74375 , n8237 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 , n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 , n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 , n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 , n8274 , n8275 , n74415 , n8277 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 , n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 , n74433 , n8295 , n8296 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 , n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n8311 , n74451 , n74452 , n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 , n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n8353 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 , n74533 , n74534 , n8396 , n8397 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 , n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 , n74553 , n74554 , n74555 , n8417 , n74557 , n74558 , n74559 , n8421 , n74561 , n74562 , n74563 , n74564 , n74565 , n8427 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 , n74573 , n74574 , n8436 , n74576 , n8438 , n8439 , n74579 , n74580 , n74581 , n74582 , n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 , n74593 , n8455 , n74595 , n74596 , n74597 , n8459 , n74599 , n74600 , n74601 , n74602 , n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 , n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 , n74633 , n74634 , n74635 , n74636 , n74637 , n8499 , n74639 , n74640 , n8502 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 , n74653 , n74654 , n74655 , n74656 , n74657 , n8519 , n8520 , n74660 , n74661 , n74662 , n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 , n74673 , n74674 , n74675 , n74676 , n74677 , n8539 , n8540 , n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 , n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n8563 , n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n8580 , n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 , n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n8602 , n8603 , n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n8619 , n74759 , n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n74776 , n74777 , n8639 , n74779 , n74780 , n74781 , n8643 , n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n8661 , n74801 , n74802 , n74803 , n8665 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 , n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n8681 , n74821 , n74822 , n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 , n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 , n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 , n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n8721 , n74861 , n74862 , n8724 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n8732 , n8733 , n74873 , n8735 , n74875 , n74876 , n74877 , n74878 , n8740 , n8741 , n74881 , n74882 , n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n8751 , n74891 , n74892 , n74893 , n74894 , n8756 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 , n74903 , n74904 , n74905 , n8767 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 , n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 , n74923 , n8785 , n74925 , n74926 , n74927 , n74928 , n74929 , n8791 , n74931 , n8793 , n8794 , n74934 , n74935 , n74936 , n8798 , n74938 , n74939 , n74940 , n8802 , n74942 , n74943 , n74944 , n8806 , n8807 , n74947 , n8809 , n74949 , n74950 , n74951 , n74952 , n8814 , n8815 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 , n74963 , n8825 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 , n74973 , n8835 , n8836 , n74976 , n74977 , n74978 , n8840 , n8841 , n74981 , n74982 , n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 , n74993 , n74994 , n74995 , n74996 , n74997 , n8859 , n8860 , n75000 , n75001 , n75002 , n75003 , n8865 , n75005 , n8867 , n8868 , n75008 , n75009 , n75010 , n8872 , n75012 , n75013 , n75014 , n8876 , n75016 , n75017 , n75018 , n8880 , n8881 , n75021 , n8883 , n75023 , n75024 , n75025 , n75026 , n8888 , n8889 , n75029 , n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n75036 , n75037 , n8899 , n75039 , n75040 , n75041 , n75042 , n8904 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 , n75053 , n8915 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 , n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n75077 , n8939 , n8940 , n75080 , n75081 , n75082 , n75083 , n8945 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 , n75093 , n8955 , n8956 , n75096 , n75097 , n75098 , n75099 , n8961 , n75101 , n8963 , n8964 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n8972 , n75112 , n75113 , n75114 , n75115 , n8977 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 , n8984 , n75124 , n75125 , n75126 , n8988 , n75128 , n75129 , n75130 , n75131 , n75132 , n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 , n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 , n9014 , n9015 , n75155 , n75156 , n75157 , n75158 , n9020 , n75160 , n75161 , n75162 , n9024 , n75164 , n75165 , n75166 , n75167 , n9029 , n9030 , n75170 , n75171 , n75172 , n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 , n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n9052 , n75192 , n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n9062 , n75202 , n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 , n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n9082 , n9083 , n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n9091 , n75231 , n75232 , n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 , n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 , n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 , n75263 , n9125 , n9126 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 , n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 , n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 , n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 , n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 , n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 , n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 , n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 , n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 , n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 , n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 , n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 , n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 , n75393 , n75394 , n9256 , n75396 , n9258 , n9259 , n75399 , n75400 , n75401 , n75402 , n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 , n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n9283 , n9284 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 , n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 , n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 , n75453 , n75454 , n75455 , n9317 , n9318 , n75458 , n75459 , n75460 , n75461 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 , n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 , n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 , n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 , n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 , n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 , n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 , n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 , n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 , n75553 , n9415 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 , n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 , n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 , n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 , n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 , n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 , n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 , n75623 , n75624 , n75625 , n9487 , n9488 , n75628 , n75629 , n75630 , n75631 , n75632 , n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 , n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 , n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 , n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 , n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 , n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 , n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 , n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 , n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 , n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 , n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 , n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 , n75753 , n75754 , n75755 , n75756 , n75757 , n9619 , n9620 , n75760 , n9622 , n9623 , n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 , n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 , n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 , n75793 , n75794 , n9656 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 , n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 , n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 , n75823 , n75824 , n75825 , n75826 , n75827 , n9689 , n75829 , n75830 , n75831 , n75832 , n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 , n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 , n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n9720 , n9721 , n75861 , n75862 , n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 , n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 , n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 , n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 , n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 , n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 , n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 , n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 , n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 , n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 , n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 , n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 , n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 , n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 , n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 , n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 , n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 , n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 , n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 , n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 , n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 , n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n9943 , n9944 , n76084 , n76085 , n76086 , n76087 , n9949 , n9950 , n76090 , n9952 , n9953 , n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 , n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 , n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n9982 , n9983 , n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 , n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 , n76143 , n76144 , n76145 , n76146 , n76147 , n10009 , n10010 , n76150 , n76151 , n76152 , n76153 , n76154 , n76155 , n76156 , n10018 , n10019 , n76159 , n76160 , n76161 , n76162 , n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 , n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 , n76183 , n76184 , n76185 , n76186 , n76187 , n10049 , n10050 , n76190 , n76191 , n76192 , n76193 , n76194 , n76195 , n76196 , n76197 , n10059 , n76199 , n76200 , n76201 , n76202 , n76203 , n76204 , n10066 , n10067 , n76207 , n10069 , n10070 , n76210 , n76211 , n76212 , n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 , n76223 , n76224 , n76225 , n76226 , n76227 , n10089 , n76229 , n76230 , n76231 , n76232 , n76233 , n76234 , n76235 , n76236 , n76237 , n10099 , n10100 , n76240 , n76241 , n76242 , n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 , n76253 , n76254 , n76255 , n76256 , n76257 , n10119 , n10120 , n76260 , n76261 , n76262 , n76263 , n76264 , n10126 , n10127 , n76267 , n10129 , n10130 , n76270 , n76271 , n76272 , n76273 , n76274 , n10136 , n10137 , n76277 , n76278 , n10140 , n76280 , n76281 , n76282 , n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 , n76293 , n76294 , n10156 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 , n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 , n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 , n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n10190 , n10191 , n76331 , n76332 , n76333 , n76334 , n10196 , n10197 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 , n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 , n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n10223 , n10224 , n76364 , n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n10232 , n10233 , n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 , n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 , n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 , n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 , n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 , n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 , n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 , n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 , n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 , n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 , n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 , n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 , n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 , n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 , n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 , n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 , n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 , n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 , n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 , n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 , n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 , n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 , n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 , n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 , n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 , n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 , n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 , n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 , n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 , n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 , n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 , n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 , n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 , n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 , n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 , n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 , n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 , n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 , n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 , n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 , n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 , n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 , n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 , n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 , n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 , n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 , n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 , n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 , n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 , n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 , n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 , n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 , n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 , n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 , n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 , n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 , n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 , n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 , n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 , n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 , n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 , n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 , n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 , n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 , n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 , n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 , n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 , n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 , n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 , n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 , n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 , n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 , n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 , n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 , n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 , n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 , n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 , n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 , n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 , n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 , n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 , n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 , n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 , n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 , n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 , n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 , n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 , n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 , n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 , n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 , n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 , n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 , n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 , n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 , n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 , n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 , n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 , n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 , n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 , n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 , n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 , n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 , n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 , n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 , n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 , n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 , n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 , n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 , n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 , n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 , n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 , n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 , n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 , n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 , n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 , n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 , n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 , n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 , n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 , n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 , n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 , n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 , n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 , n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 , n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 , n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 , n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 , n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 , n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 , n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 , n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 , n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 , n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 , n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 , n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 , n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 , n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 , n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 , n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 , n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 , n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782;
buf ( n243 , n2533 );
buf ( n244 , n2538 );
buf ( n245 , n2543 );
buf ( n246 , n2548 );
buf ( n247 , n2553 );
buf ( n248 , n2558 );
buf ( n249 , n2563 );
buf ( n250 , n2568 );
buf ( n251 , n2573 );
buf ( n252 , n2578 );
buf ( n253 , n2583 );
buf ( n254 , n2588 );
buf ( n255 , n2593 );
buf ( n256 , n2598 );
buf ( n257 , n2603 );
buf ( n258 , n2605 );
buf ( n259 , n68749 );
buf ( n260 , n68751 );
buf ( n261 , n68756 );
buf ( n262 , n2622 );
buf ( n263 , n2624 );
buf ( n264 , n68765 );
buf ( n265 , n2628 );
buf ( n266 , n68769 );
buf ( n267 , n68771 );
buf ( n268 , n2634 );
buf ( n269 , n2636 );
buf ( n270 , n2638 );
buf ( n271 , n68779 );
buf ( n272 , n68781 );
buf ( n273 , n2644 );
buf ( n274 , n68785 );
buf ( n275 , n2648 );
buf ( n276 , n2650 );
buf ( n277 , n2652 );
buf ( n278 , n2654 );
buf ( n279 , n68795 );
buf ( n280 , n2658 );
buf ( n281 , n68799 );
buf ( n282 , n68801 );
buf ( n283 , n2664 );
buf ( n284 , n2666 );
buf ( n285 , n2668 );
buf ( n286 , n68809 );
buf ( n287 , n68811 );
buf ( n288 , n2674 );
buf ( n289 , n68815 );
buf ( n290 , n2681 );
buf ( n291 , n68825 );
buf ( n292 , n2688 );
buf ( n293 , n68829 );
buf ( n294 , n68831 );
buf ( PO_rd , n2694 );
buf ( PO_wr , n2696 );
buf ( DFF_state_reg_S , n71972 );
buf ( DFF_state_reg_R , n71974 );
buf ( DFF_state_reg_CK , n71975 );
buf ( DFF_state_reg_D , n71976 );
buf ( n295 , n76381 );
buf ( n296 , n76383 );
buf ( n297 , n76384 );
buf ( n298 , n76390 );
buf ( n299 , n10137 );
buf ( n300 , n76278 );
buf ( n301 , n10140 );
buf ( n302 , n76285 );
buf ( n303 , n76167 );
buf ( n304 , n76169 );
buf ( n305 , n76170 );
buf ( n306 , n76176 );
buf ( n307 , n76139 );
buf ( n308 , n76141 );
buf ( n309 , n76142 );
buf ( n310 , n10009 );
buf ( n311 , n76129 );
buf ( n312 , n76131 );
buf ( n313 , n76132 );
buf ( n314 , n76138 );
buf ( n315 , n76119 );
buf ( n316 , n9982 );
buf ( n317 , n9983 );
buf ( n318 , n76128 );
buf ( n319 , n76109 );
buf ( n320 , n76111 );
buf ( n321 , n76112 );
buf ( n322 , n76118 );
buf ( n323 , n76099 );
buf ( n324 , n76101 );
buf ( n325 , n76102 );
buf ( n326 , n76108 );
buf ( n327 , n9950 );
buf ( n328 , n9952 );
buf ( n329 , n9953 );
buf ( n330 , n76098 );
buf ( n331 , n76080 );
buf ( n332 , n9943 );
buf ( n333 , n9944 );
buf ( n334 , n9949 );
buf ( n335 , n10233 );
buf ( n336 , n76374 );
buf ( n337 , n76375 );
buf ( n338 , n76380 );
buf ( n339 , n10224 );
buf ( n340 , n76365 );
buf ( n341 , n76366 );
buf ( n342 , n10232 );
buf ( n343 , n76354 );
buf ( n344 , n76356 );
buf ( n345 , n76357 );
buf ( n346 , n10223 );
buf ( n347 , n76345 );
buf ( n348 , n76347 );
buf ( n349 , n76348 );
buf ( n350 , n76353 );
buf ( n351 , n10197 );
buf ( n352 , n76338 );
buf ( n353 , n76339 );
buf ( n354 , n76344 );
buf ( n355 , n76327 );
buf ( n356 , n10190 );
buf ( n357 , n10191 );
buf ( n358 , n10196 );
buf ( n359 , n76317 );
buf ( n360 , n76319 );
buf ( n361 , n76320 );
buf ( n362 , n76326 );
buf ( n363 , n76307 );
buf ( n364 , n76309 );
buf ( n365 , n76310 );
buf ( n366 , n76316 );
buf ( n367 , n76296 );
buf ( n368 , n76298 );
buf ( n369 , n76299 );
buf ( n370 , n76306 );
buf ( n371 , n76286 );
buf ( n372 , n76288 );
buf ( n373 , n76289 );
buf ( n374 , n10156 );
buf ( n375 , n10127 );
buf ( n376 , n10129 );
buf ( n377 , n10130 );
buf ( n378 , n10136 );
buf ( n379 , n76256 );
buf ( n380 , n10119 );
buf ( n381 , n10120 );
buf ( n382 , n10126 );
buf ( n383 , n76246 );
buf ( n384 , n76248 );
buf ( n385 , n76249 );
buf ( n386 , n76255 );
buf ( n387 , n76236 );
buf ( n388 , n10099 );
buf ( n389 , n10100 );
buf ( n390 , n76245 );
buf ( n391 , n76226 );
buf ( n392 , n10089 );
buf ( n393 , n76229 );
buf ( n394 , n76235 );
buf ( n395 , n76216 );
buf ( n396 , n76218 );
buf ( n397 , n76219 );
buf ( n398 , n76225 );
buf ( n399 , n10067 );
buf ( n400 , n10069 );
buf ( n401 , n10070 );
buf ( n402 , n76215 );
buf ( n403 , n76196 );
buf ( n404 , n10059 );
buf ( n405 , n76199 );
buf ( n406 , n10066 );
buf ( n407 , n76186 );
buf ( n408 , n10049 );
buf ( n409 , n10050 );
buf ( n410 , n76195 );
buf ( n411 , n76177 );
buf ( n412 , n76179 );
buf ( n413 , n76180 );
buf ( n414 , n76185 );
buf ( n415 , n10019 );
buf ( n416 , n76160 );
buf ( n417 , n76161 );
buf ( n418 , n76166 );
buf ( n419 , n10010 );
buf ( n420 , n76151 );
buf ( n421 , n76152 );
buf ( n422 , n10018 );
buf ( n423 , n75253 );
buf ( n424 , n75255 );
buf ( n425 , n75256 );
buf ( n426 , n75261 );
buf ( n427 , n75243 );
buf ( n428 , n75245 );
buf ( n429 , n75246 );
buf ( n430 , n75252 );
buf ( n431 , n73725 );
buf ( n432 , n73727 );
buf ( n433 , n73728 );
buf ( n434 , n7619 );
buf ( n435 , n73404 );
buf ( n436 , n73406 );
buf ( n437 , n73407 );
buf ( n438 , n73440 );
buf ( n439 , n72376 );
buf ( n440 , n72378 );
buf ( n441 , n72379 );
buf ( n442 , n72424 );
buf ( n443 , n6185 );
buf ( n444 , n72326 );
buf ( n445 , n72327 );
buf ( n446 , n72375 );
buf ( n447 , n6137 );
buf ( n448 , n72278 );
buf ( n449 , n72279 );
buf ( n450 , n6184 );
buf ( n451 , n72214 );
buf ( n452 , n6077 );
buf ( n453 , n72217 );
buf ( n454 , n6136 );
buf ( n455 , n72157 );
buf ( n456 , n72159 );
buf ( n457 , n6021 );
buf ( n458 , n72213 );
buf ( n459 , n72078 );
buf ( n460 , n72080 );
buf ( n461 , n72081 );
buf ( n462 , n6017 );
buf ( n463 , n72026 );
buf ( n464 , n5889 );
buf ( n465 , n72029 );
buf ( n466 , n72077 );
buf ( n467 , n71977 );
buf ( n468 , n71979 );
buf ( n469 , n71980 );
buf ( n470 , n72025 );
buf ( n471 , n73700 );
buf ( n472 , n73702 );
buf ( n473 , n73703 );
buf ( n474 , n73724 );
buf ( n475 , n7537 );
buf ( n476 , n7539 );
buf ( n477 , n7540 );
buf ( n478 , n73699 );
buf ( n479 , n73651 );
buf ( n480 , n73653 );
buf ( n481 , n73654 );
buf ( n482 , n7536 );
buf ( n483 , n73577 );
buf ( n484 , n73579 );
buf ( n485 , n73580 );
buf ( n486 , n73650 );
buf ( n487 , n73553 );
buf ( n488 , n73555 );
buf ( n489 , n73556 );
buf ( n490 , n73576 );
buf ( n491 , n7389 );
buf ( n492 , n7391 );
buf ( n493 , n7392 );
buf ( n494 , n73552 );
buf ( n495 , n73508 );
buf ( n496 , n73510 );
buf ( n497 , n73511 );
buf ( n498 , n7388 );
buf ( n499 , n73486 );
buf ( n500 , n7349 );
buf ( n501 , n7350 );
buf ( n502 , n73507 );
buf ( n503 , n73464 );
buf ( n504 , n7327 );
buf ( n505 , n7328 );
buf ( n506 , n73485 );
buf ( n507 , n73441 );
buf ( n508 , n73443 );
buf ( n509 , n7305 );
buf ( n510 , n73463 );
buf ( n511 , n7208 );
buf ( n512 , n73349 );
buf ( n513 , n73350 );
buf ( n514 , n73403 );
buf ( n515 , n73276 );
buf ( n516 , n7139 );
buf ( n517 , n73279 );
buf ( n518 , n7207 );
buf ( n519 , n73212 );
buf ( n520 , n73214 );
buf ( n521 , n73215 );
buf ( n522 , n73275 );
buf ( n523 , n73127 );
buf ( n524 , n73129 );
buf ( n525 , n6991 );
buf ( n526 , n73211 );
buf ( n527 , n6927 );
buf ( n528 , n73068 );
buf ( n529 , n73069 );
buf ( n530 , n6987 );
buf ( n531 , n72992 );
buf ( n532 , n72994 );
buf ( n533 , n6856 );
buf ( n534 , n6926 );
buf ( n535 , n6777 );
buf ( n536 , n72918 );
buf ( n537 , n72919 );
buf ( n538 , n6852 );
buf ( n539 , n72833 );
buf ( n540 , n6696 );
buf ( n541 , n72836 );
buf ( n542 , n6776 );
buf ( n543 , n72425 );
buf ( n544 , n72427 );
buf ( n545 , n72428 );
buf ( n546 , n72832 );
buf ( n547 , n74841 );
buf ( n548 , n74843 );
buf ( n549 , n74844 );
buf ( n550 , n8721 );
buf ( n551 , n74801 );
buf ( n552 , n74803 );
buf ( n553 , n8665 );
buf ( n554 , n74819 );
buf ( n555 , n8436 );
buf ( n556 , n8438 );
buf ( n557 , n8439 );
buf ( n558 , n8455 );
buf ( n559 , n8397 );
buf ( n560 , n74538 );
buf ( n561 , n74539 );
buf ( n562 , n8417 );
buf ( n563 , n74514 );
buf ( n564 , n74516 );
buf ( n565 , n74517 );
buf ( n566 , n8396 );
buf ( n567 , n8353 );
buf ( n568 , n74494 );
buf ( n569 , n74495 );
buf ( n570 , n74513 );
buf ( n571 , n74474 );
buf ( n572 , n74476 );
buf ( n573 , n74477 );
buf ( n574 , n74491 );
buf ( n575 , n8311 );
buf ( n576 , n74452 );
buf ( n577 , n74453 );
buf ( n578 , n74473 );
buf ( n579 , n74432 );
buf ( n580 , n8295 );
buf ( n581 , n8296 );
buf ( n582 , n74449 );
buf ( n583 , n70906 );
buf ( n584 , n4769 );
buf ( n585 , n4770 );
buf ( n586 , n4881 );
buf ( n587 , n71659 );
buf ( n588 , n71661 );
buf ( n589 , n71662 );
buf ( n590 , n71718 );
buf ( n591 , n5440 );
buf ( n592 , n71581 );
buf ( n593 , n71582 );
buf ( n594 , n71658 );
buf ( n595 , n5374 );
buf ( n596 , n71515 );
buf ( n597 , n71516 );
buf ( n598 , n5439 );
buf ( n599 , n8681 );
buf ( n600 , n74822 );
buf ( n601 , n74823 );
buf ( n602 , n74840 );
buf ( n603 , n71440 );
buf ( n604 , n71442 );
buf ( n605 , n5304 );
buf ( n606 , n71512 );
buf ( n607 , n71348 );
buf ( n608 , n71350 );
buf ( n609 , n71351 );
buf ( n610 , n5300 );
buf ( n611 , n71324 );
buf ( n612 , n71326 );
buf ( n613 , n71327 );
buf ( n614 , n71347 );
buf ( n615 , n71268 );
buf ( n616 , n71270 );
buf ( n617 , n5132 );
buf ( n618 , n71323 );
buf ( n619 , n5072 );
buf ( n620 , n5074 );
buf ( n621 , n5075 );
buf ( n622 , n5128 );
buf ( n623 , n71021 );
buf ( n624 , n4884 );
buf ( n625 , n4885 );
buf ( n626 , n5071 );
buf ( n627 , n74779 );
buf ( n628 , n74781 );
buf ( n629 , n8643 );
buf ( n630 , n8661 );
buf ( n631 , n74759 );
buf ( n632 , n74761 );
buf ( n633 , n74762 );
buf ( n634 , n8639 );
buf ( n635 , n74739 );
buf ( n636 , n8602 );
buf ( n637 , n8603 );
buf ( n638 , n8619 );
buf ( n639 , n8580 );
buf ( n640 , n74721 );
buf ( n641 , n74722 );
buf ( n642 , n74738 );
buf ( n643 , n74699 );
buf ( n644 , n74701 );
buf ( n645 , n8563 );
buf ( n646 , n74718 );
buf ( n647 , n8540 );
buf ( n648 , n74681 );
buf ( n649 , n74682 );
buf ( n650 , n74698 );
buf ( n651 , n8520 );
buf ( n652 , n74661 );
buf ( n653 , n74662 );
buf ( n654 , n8539 );
buf ( n655 , n74639 );
buf ( n656 , n8502 );
buf ( n657 , n74642 );
buf ( n658 , n8519 );
buf ( n659 , n74617 );
buf ( n660 , n74619 );
buf ( n661 , n74620 );
buf ( n662 , n8499 );
buf ( n663 , n74595 );
buf ( n664 , n74597 );
buf ( n665 , n8459 );
buf ( n666 , n74616 );
buf ( n667 , n8427 );
buf ( n668 , n74568 );
buf ( n669 , n74569 );
buf ( n670 , n74574 );
buf ( n671 , n74557 );
buf ( n672 , n74559 );
buf ( n673 , n8421 );
buf ( n674 , n74565 );
buf ( n675 , n8977 );
buf ( n676 , n75118 );
buf ( n677 , n75119 );
buf ( n678 , n8984 );
buf ( n679 , n8889 );
buf ( n680 , n75030 );
buf ( n681 , n75031 );
buf ( n682 , n75035 );
buf ( n683 , n74938 );
buf ( n684 , n74940 );
buf ( n685 , n8802 );
buf ( n686 , n8806 );
buf ( n687 , n74912 );
buf ( n688 , n74914 );
buf ( n689 , n74915 );
buf ( n690 , n74920 );
buf ( n691 , n74904 );
buf ( n692 , n8767 );
buf ( n693 , n74907 );
buf ( n694 , n74911 );
buf ( n695 , n74896 );
buf ( n696 , n74898 );
buf ( n697 , n74899 );
buf ( n698 , n74903 );
buf ( n699 , n74888 );
buf ( n700 , n8751 );
buf ( n701 , n74891 );
buf ( n702 , n8756 );
buf ( n703 , n8741 );
buf ( n704 , n74882 );
buf ( n705 , n74883 );
buf ( n706 , n74887 );
buf ( n707 , n8733 );
buf ( n708 , n8735 );
buf ( n709 , n74875 );
buf ( n710 , n8740 );
buf ( n711 , n74861 );
buf ( n712 , n8724 );
buf ( n713 , n74864 );
buf ( n714 , n8732 );
buf ( n715 , n75108 );
buf ( n716 , n75110 );
buf ( n717 , n8972 );
buf ( n718 , n75115 );
buf ( n719 , n8961 );
buf ( n720 , n8963 );
buf ( n721 , n8964 );
buf ( n722 , n75107 );
buf ( n723 , n75092 );
buf ( n724 , n8955 );
buf ( n725 , n8956 );
buf ( n726 , n75099 );
buf ( n727 , n8945 );
buf ( n728 , n75086 );
buf ( n729 , n75087 );
buf ( n730 , n75091 );
buf ( n731 , n75076 );
buf ( n732 , n8939 );
buf ( n733 , n8940 );
buf ( n734 , n75083 );
buf ( n735 , n75068 );
buf ( n736 , n75070 );
buf ( n737 , n75071 );
buf ( n738 , n75075 );
buf ( n739 , n75060 );
buf ( n740 , n75062 );
buf ( n741 , n75063 );
buf ( n742 , n75067 );
buf ( n743 , n75052 );
buf ( n744 , n8915 );
buf ( n745 , n75055 );
buf ( n746 , n75059 );
buf ( n747 , n75044 );
buf ( n748 , n75046 );
buf ( n749 , n75047 );
buf ( n750 , n75051 );
buf ( n751 , n75036 );
buf ( n752 , n8899 );
buf ( n753 , n75039 );
buf ( n754 , n8904 );
buf ( n755 , n8881 );
buf ( n756 , n8883 );
buf ( n757 , n75023 );
buf ( n758 , n8888 );
buf ( n759 , n75012 );
buf ( n760 , n75014 );
buf ( n761 , n8876 );
buf ( n762 , n8880 );
buf ( n763 , n8865 );
buf ( n764 , n8867 );
buf ( n765 , n8868 );
buf ( n766 , n8872 );
buf ( n767 , n74996 );
buf ( n768 , n8859 );
buf ( n769 , n8860 );
buf ( n770 , n75003 );
buf ( n771 , n74988 );
buf ( n772 , n74990 );
buf ( n773 , n74991 );
buf ( n774 , n74995 );
buf ( n775 , n8841 );
buf ( n776 , n74982 );
buf ( n777 , n74983 );
buf ( n778 , n74987 );
buf ( n779 , n74972 );
buf ( n780 , n8835 );
buf ( n781 , n8836 );
buf ( n782 , n8840 );
buf ( n783 , n74962 );
buf ( n784 , n8825 );
buf ( n785 , n74965 );
buf ( n786 , n74971 );
buf ( n787 , n8815 );
buf ( n788 , n74956 );
buf ( n789 , n74957 );
buf ( n790 , n74961 );
buf ( n791 , n8807 );
buf ( n792 , n8809 );
buf ( n793 , n74949 );
buf ( n794 , n8814 );
buf ( n795 , n8791 );
buf ( n796 , n8793 );
buf ( n797 , n8794 );
buf ( n798 , n8798 );
buf ( n799 , n74921 );
buf ( n800 , n74923 );
buf ( n801 , n8785 );
buf ( n802 , n74929 );
buf ( DFF_B_reg_S , n76391 );
buf ( DFF_B_reg_R , n76393 );
buf ( DFF_B_reg_CK , n76394 );
buf ( DFF_B_reg_D , n77765 );
buf ( n803 , n8275 );
buf ( n804 , n8277 );
buf ( n805 , n74417 );
buf ( n806 , n74431 );
buf ( n807 , n8084 );
buf ( n808 , n74225 );
buf ( n809 , n74226 );
buf ( n810 , n74243 );
buf ( n811 , n73952 );
buf ( n812 , n73954 );
buf ( n813 , n73955 );
buf ( n814 , n7829 );
buf ( n815 , n73873 );
buf ( n816 , n73875 );
buf ( n817 , n73876 );
buf ( n818 , n7749 );
buf ( n819 , n73850 );
buf ( n820 , n73852 );
buf ( n821 , n7714 );
buf ( n822 , n73872 );
buf ( n823 , n7693 );
buf ( n824 , n73834 );
buf ( n825 , n7696 );
buf ( n826 , n73849 );
buf ( n827 , n7677 );
buf ( n828 , n73818 );
buf ( n829 , n73819 );
buf ( n830 , n7692 );
buf ( n831 , n73800 );
buf ( n832 , n73802 );
buf ( n833 , n73803 );
buf ( n834 , n7676 );
buf ( n835 , n7641 );
buf ( n836 , n73782 );
buf ( n837 , n73783 );
buf ( n838 , n73799 );
buf ( n839 , n73759 );
buf ( n840 , n7622 );
buf ( n841 , n7623 );
buf ( n842 , n7640 );
buf ( n843 , n74395 );
buf ( n844 , n74397 );
buf ( n845 , n74398 );
buf ( n846 , n8274 );
buf ( n847 , n8237 );
buf ( n848 , n74378 );
buf ( n849 , n74379 );
buf ( n850 , n74394 );
buf ( n851 , n74357 );
buf ( n852 , n74359 );
buf ( n853 , n8221 );
buf ( n854 , n74375 );
buf ( n855 , n8199 );
buf ( n856 , n8201 );
buf ( n857 , n8202 );
buf ( n858 , n8217 );
buf ( n859 , n74319 );
buf ( n860 , n74321 );
buf ( n861 , n74322 );
buf ( n862 , n74337 );
buf ( n863 , n74300 );
buf ( n864 , n8163 );
buf ( n865 , n8164 );
buf ( n866 , n74318 );
buf ( n867 , n2698 );
buf ( n868 , n68840 );
buf ( n869 , n68841 );
buf ( n870 , n70905 );
buf ( n871 , n8143 );
buf ( n872 , n74284 );
buf ( n873 , n74285 );
buf ( n874 , n74299 );
buf ( n875 , n74263 );
buf ( n876 , n8126 );
buf ( n877 , n8127 );
buf ( n878 , n8142 );
buf ( n879 , n74244 );
buf ( n880 , n74246 );
buf ( n881 , n74247 );
buf ( n882 , n74262 );
buf ( n883 , n74204 );
buf ( n884 , n8067 );
buf ( n885 , n8068 );
buf ( n886 , n74222 );
buf ( n887 , n8046 );
buf ( n888 , n74187 );
buf ( n889 , n74188 );
buf ( n890 , n74203 );
buf ( n891 , n8027 );
buf ( n892 , n74168 );
buf ( n893 , n74169 );
buf ( n894 , n8045 );
buf ( n895 , n74147 );
buf ( n896 , n8010 );
buf ( n897 , n8011 );
buf ( n898 , n8026 );
buf ( n899 , n7989 );
buf ( n900 , n74130 );
buf ( n901 , n7992 );
buf ( n902 , n74146 );
buf ( n903 , n7972 );
buf ( n904 , n74113 );
buf ( n905 , n74114 );
buf ( n906 , n7988 );
buf ( n907 , n74093 );
buf ( n908 , n74095 );
buf ( n909 , n74096 );
buf ( n910 , n7971 );
buf ( n911 , n7937 );
buf ( n912 , n74078 );
buf ( n913 , n74079 );
buf ( n914 , n7953 );
buf ( n915 , n7921 );
buf ( n916 , n74062 );
buf ( n917 , n74063 );
buf ( n918 , n7936 );
buf ( n919 , n7830 );
buf ( n920 , n7832 );
buf ( n921 , n7833 );
buf ( n922 , n7920 );
buf ( n923 , n7793 );
buf ( n924 , n73934 );
buf ( n925 , n73935 );
buf ( n926 , n73951 );
buf ( n927 , n7750 );
buf ( n928 , n73891 );
buf ( n929 , n73892 );
buf ( n930 , n73931 );
buf ( n931 , n76066 );
buf ( n932 , n76068 );
buf ( n933 , n76069 );
buf ( n934 , n76079 );
buf ( n935 , n75608 );
buf ( n936 , n75610 );
buf ( n937 , n75611 );
buf ( n938 , n75623 );
buf ( n939 , n75578 );
buf ( n940 , n75580 );
buf ( n941 , n75581 );
buf ( n942 , n75607 );
buf ( n943 , n75551 );
buf ( n944 , n75553 );
buf ( n945 , n9415 );
buf ( n946 , n75577 );
buf ( n947 , n75515 );
buf ( n948 , n75517 );
buf ( n949 , n75518 );
buf ( n950 , n75550 );
buf ( n951 , n75484 );
buf ( n952 , n75486 );
buf ( n953 , n75487 );
buf ( n954 , n75514 );
buf ( n955 , n9318 );
buf ( n956 , n75459 );
buf ( n957 , n75460 );
buf ( n958 , n75483 );
buf ( n959 , n75420 );
buf ( n960 , n9283 );
buf ( n961 , n9284 );
buf ( n962 , n9317 );
buf ( n963 , n9256 );
buf ( n964 , n9258 );
buf ( n965 , n9259 );
buf ( n966 , n75419 );
buf ( n967 , n75262 );
buf ( n968 , n9125 );
buf ( n969 , n9126 );
buf ( n970 , n75394 );
buf ( n971 , n76038 );
buf ( n972 , n76040 );
buf ( n973 , n76041 );
buf ( n974 , n76065 );
buf ( n975 , n76000 );
buf ( n976 , n76002 );
buf ( n977 , n76003 );
buf ( n978 , n76037 );
buf ( n979 , n75974 );
buf ( n980 , n75976 );
buf ( n981 , n75977 );
buf ( n982 , n75999 );
buf ( n983 , n75940 );
buf ( n984 , n75942 );
buf ( n985 , n75943 );
buf ( n986 , n75973 );
buf ( n987 , n75910 );
buf ( n988 , n75912 );
buf ( n989 , n75913 );
buf ( n990 , n75939 );
buf ( n991 , n9721 );
buf ( n992 , n75862 );
buf ( n993 , n75863 );
buf ( n994 , n75909 );
buf ( n995 , n75829 );
buf ( n996 , n75831 );
buf ( n997 , n75832 );
buf ( n998 , n9720 );
buf ( n999 , n75796 );
buf ( n1000 , n75798 );
buf ( n1001 , n75799 );
buf ( n1002 , n9689 );
buf ( n1003 , n9620 );
buf ( n1004 , n9622 );
buf ( n1005 , n9623 );
buf ( n1006 , n9656 );
buf ( n1007 , n75624 );
buf ( n1008 , n9487 );
buf ( n1009 , n9488 );
buf ( n1010 , n9619 );
buf ( n1011 , n75231 );
buf ( n1012 , n75233 );
buf ( n1013 , n75234 );
buf ( n1014 , n75242 );
buf ( n1015 , n75219 );
buf ( n1016 , n9082 );
buf ( n1017 , n9083 );
buf ( n1018 , n9091 );
buf ( n1019 , n75189 );
buf ( n1020 , n9052 );
buf ( n1021 , n75192 );
buf ( n1022 , n75200 );
buf ( n1023 , n9030 );
buf ( n1024 , n75171 );
buf ( n1025 , n75172 );
buf ( n1026 , n75179 );
buf ( n1027 , n75160 );
buf ( n1028 , n75162 );
buf ( n1029 , n9024 );
buf ( n1030 , n9029 );
buf ( n1031 , n75151 );
buf ( n1032 , n9014 );
buf ( n1033 , n9015 );
buf ( n1034 , n9020 );
buf ( n1035 , n75142 );
buf ( n1036 , n75144 );
buf ( n1037 , n75145 );
buf ( n1038 , n75150 );
buf ( n1039 , n75133 );
buf ( n1040 , n75135 );
buf ( n1041 , n75136 );
buf ( n1042 , n75141 );
buf ( n1043 , n75124 );
buf ( n1044 , n75126 );
buf ( n1045 , n8988 );
buf ( n1046 , n75132 );
buf ( n1047 , n71719 );
buf ( n1048 , n5582 );
buf ( n1049 , n71722 );
buf ( n1050 , n5591 );
buf ( n1051 , n71963 );
buf ( n1052 , n71965 );
buf ( n1053 , n71966 );
buf ( n1054 , n71971 );
buf ( n1055 , n71954 );
buf ( n1056 , n71956 );
buf ( n1057 , n71957 );
buf ( n1058 , n71962 );
buf ( n1059 , n71945 );
buf ( n1060 , n71947 );
buf ( n1061 , n71948 );
buf ( n1062 , n71953 );
buf ( n1063 , n71936 );
buf ( n1064 , n71938 );
buf ( n1065 , n71939 );
buf ( n1066 , n71944 );
buf ( n1067 , n71927 );
buf ( n1068 , n71929 );
buf ( n1069 , n71930 );
buf ( n1070 , n71935 );
buf ( n1071 , n71918 );
buf ( n1072 , n71920 );
buf ( n1073 , n71921 );
buf ( n1074 , n71926 );
buf ( n1075 , n71909 );
buf ( n1076 , n71911 );
buf ( n1077 , n71912 );
buf ( n1078 , n71917 );
buf ( n1079 , n71900 );
buf ( n1080 , n71902 );
buf ( n1081 , n71903 );
buf ( n1082 , n71908 );
buf ( n1083 , n5752 );
buf ( n1084 , n5754 );
buf ( n1085 , n5755 );
buf ( n1086 , n71899 );
buf ( n1087 , n71882 );
buf ( n1088 , n5745 );
buf ( n1089 , n71885 );
buf ( n1090 , n5751 );
buf ( n1091 , n5734 );
buf ( n1092 , n71875 );
buf ( n1093 , n71876 );
buf ( n1094 , n5742 );
buf ( n1095 , n71856 );
buf ( n1096 , n71858 );
buf ( n1097 , n71859 );
buf ( n1098 , n71872 );
buf ( n1099 , n71838 );
buf ( n1100 , n5701 );
buf ( n1101 , n5702 );
buf ( n1102 , n71855 );
buf ( n1103 , n71818 );
buf ( n1104 , n5681 );
buf ( n1105 , n5682 );
buf ( n1106 , n71837 );
buf ( n1107 , n5664 );
buf ( n1108 , n71805 );
buf ( n1109 , n71806 );
buf ( n1110 , n71817 );
buf ( n1111 , n5645 );
buf ( n1112 , n71786 );
buf ( n1113 , n71787 );
buf ( n1114 , n71802 );
buf ( n1115 , n71767 );
buf ( n1116 , n71769 );
buf ( n1117 , n5631 );
buf ( n1118 , n5644 );
buf ( n1119 , n5601 );
buf ( n1120 , n71742 );
buf ( n1121 , n5604 );
buf ( n1122 , n71766 );
buf ( n1123 , n75210 );
buf ( n1124 , n75212 );
buf ( n1125 , n75213 );
buf ( n1126 , n75218 );
buf ( n1127 , n9062 );
buf ( n1128 , n75203 );
buf ( n1129 , n75204 );
buf ( n1130 , n75209 );
buf ( n1131 , n75180 );
buf ( n1132 , n75182 );
buf ( n1133 , n75183 );
buf ( n1134 , n75188 );
buf ( n1135 , n5592 );
buf ( n1136 , n5594 );
buf ( n1137 , n5595 );
buf ( n1138 , n71739 );
buf ( DFF_rd_reg_S , n77772 );
buf ( DFF_rd_reg_R , n77774 );
buf ( DFF_rd_reg_CK , n77775 );
buf ( DFF_rd_reg_D , n77782 );
buf ( DFF_wr_reg_S , n77766 );
buf ( DFF_wr_reg_R , n77769 );
buf ( DFF_wr_reg_CK , n77770 );
buf ( DFF_wr_reg_D , n77771 );
buf ( n68634 , PI_clock );
buf ( n68635 , PI_reset );
buf ( n68636 , n0 );
buf ( n2498 , n1 );
buf ( n2499 , n2 );
buf ( n2500 , n3 );
buf ( n2501 , n4 );
buf ( n2502 , n5 );
buf ( n2503 , n6 );
buf ( n2504 , n7 );
buf ( n68644 , n8 );
buf ( n68645 , n9 );
buf ( n68646 , n10 );
buf ( n2508 , n11 );
buf ( n2509 , n12 );
buf ( n68649 , n13 );
buf ( n68650 , n14 );
buf ( n68651 , n15 );
buf ( n2513 , n16 );
buf ( n2514 , n17 );
buf ( n2515 , n18 );
buf ( n2516 , n19 );
buf ( n2517 , n20 );
buf ( n2518 , n21 );
buf ( n2519 , n22 );
buf ( n68659 , n23 );
buf ( n68660 , n24 );
buf ( n68661 , n25 );
buf ( n2523 , n26 );
buf ( n2524 , n27 );
buf ( n68664 , n28 );
buf ( n68665 , n29 );
buf ( n68666 , n30 );
buf ( n2528 , n31 );
buf ( n2529 , n210 );
not ( n68669 , n2529 );
not ( n68670 , n68669 );
buf ( n2532 , n68670 );
buf ( n2533 , n2532 );
buf ( n2534 , n209 );
not ( n68674 , n2534 );
not ( n68675 , n68674 );
buf ( n68676 , n68675 );
buf ( n2538 , n68676 );
buf ( n2539 , n208 );
not ( n68679 , n2539 );
not ( n68680 , n68679 );
buf ( n68681 , n68680 );
buf ( n2543 , n68681 );
buf ( n2544 , n207 );
not ( n68684 , n2544 );
not ( n68685 , n68684 );
buf ( n2547 , n68685 );
buf ( n2548 , n2547 );
buf ( n2549 , n206 );
not ( n68689 , n2549 );
not ( n68690 , n68689 );
buf ( n68691 , n68690 );
buf ( n2553 , n68691 );
buf ( n2554 , n205 );
not ( n68694 , n2554 );
not ( n68695 , n68694 );
buf ( n68696 , n68695 );
buf ( n2558 , n68696 );
buf ( n2559 , n204 );
not ( n68699 , n2559 );
not ( n68700 , n68699 );
buf ( n2562 , n68700 );
buf ( n2563 , n2562 );
buf ( n2564 , n203 );
not ( n68704 , n2564 );
not ( n68705 , n68704 );
buf ( n68706 , n68705 );
buf ( n2568 , n68706 );
buf ( n2569 , n202 );
not ( n68709 , n2569 );
not ( n68710 , n68709 );
buf ( n68711 , n68710 );
buf ( n2573 , n68711 );
buf ( n2574 , n201 );
not ( n68714 , n2574 );
not ( n68715 , n68714 );
buf ( n2577 , n68715 );
buf ( n2578 , n2577 );
buf ( n2579 , n200 );
not ( n68719 , n2579 );
not ( n68720 , n68719 );
buf ( n68721 , n68720 );
buf ( n2583 , n68721 );
buf ( n2584 , n199 );
not ( n68724 , n2584 );
not ( n68725 , n68724 );
buf ( n68726 , n68725 );
buf ( n2588 , n68726 );
buf ( n2589 , n198 );
not ( n68729 , n2589 );
not ( n68730 , n68729 );
buf ( n2592 , n68730 );
buf ( n2593 , n2592 );
buf ( n2594 , n197 );
not ( n68734 , n2594 );
not ( n68735 , n68734 );
buf ( n68736 , n68735 );
buf ( n2598 , n68736 );
buf ( n2599 , n196 );
not ( n68739 , n2599 );
not ( n68740 , n68739 );
buf ( n68741 , n68740 );
buf ( n2603 , n68741 );
buf ( n2604 , n195 );
buf ( n2605 , n2604 );
buf ( n2606 , n194 );
not ( n68746 , n2606 );
not ( n68747 , n68746 );
buf ( n2609 , n68747 );
buf ( n68749 , n2609 );
buf ( n68750 , n193 );
buf ( n68751 , n68750 );
buf ( n2613 , n192 );
not ( n68753 , n2613 );
not ( n68754 , n68753 );
buf ( n68755 , n68754 );
buf ( n68756 , n68755 );
buf ( n2618 , n191 );
not ( n68758 , n2618 );
not ( n68759 , n68758 );
buf ( n2621 , n68759 );
buf ( n2622 , n2621 );
buf ( n2623 , n242 );
buf ( n2624 , n2623 );
buf ( n68764 , n241 );
buf ( n68765 , n68764 );
buf ( n68766 , n240 );
buf ( n2628 , n68766 );
buf ( n2629 , n239 );
buf ( n68769 , n2629 );
buf ( n68770 , n238 );
buf ( n68771 , n68770 );
buf ( n2633 , n237 );
buf ( n2634 , n2633 );
buf ( n2635 , n236 );
buf ( n2636 , n2635 );
buf ( n2637 , n235 );
buf ( n2638 , n2637 );
buf ( n2639 , n234 );
buf ( n68779 , n2639 );
buf ( n68780 , n233 );
buf ( n68781 , n68780 );
buf ( n2643 , n232 );
buf ( n2644 , n2643 );
buf ( n68784 , n231 );
buf ( n68785 , n68784 );
buf ( n68786 , n230 );
buf ( n2648 , n68786 );
buf ( n2649 , n229 );
buf ( n2650 , n2649 );
buf ( n2651 , n228 );
buf ( n2652 , n2651 );
buf ( n2653 , n227 );
buf ( n2654 , n2653 );
buf ( n68794 , n226 );
buf ( n68795 , n68794 );
buf ( n68796 , n225 );
buf ( n2658 , n68796 );
buf ( n2659 , n224 );
buf ( n68799 , n2659 );
buf ( n68800 , n223 );
buf ( n68801 , n68800 );
buf ( n2663 , n222 );
buf ( n2664 , n2663 );
buf ( n2665 , n221 );
buf ( n2666 , n2665 );
buf ( n2667 , n220 );
buf ( n2668 , n2667 );
buf ( n2669 , n219 );
buf ( n68809 , n2669 );
buf ( n68810 , n218 );
buf ( n68811 , n68810 );
buf ( n2673 , n217 );
buf ( n2674 , n2673 );
buf ( n68814 , n216 );
buf ( n68815 , n68814 );
buf ( n68816 , n215 );
not ( n68817 , n68816 );
not ( n68818 , n68817 );
buf ( n2680 , n68818 );
buf ( n2681 , n2680 );
buf ( n2682 , n214 );
not ( n68822 , n2682 );
not ( n68823 , n68822 );
buf ( n68824 , n68823 );
buf ( n68825 , n68824 );
buf ( n68826 , n213 );
buf ( n2688 , n68826 );
buf ( n2689 , n212 );
buf ( n68829 , n2689 );
buf ( n68830 , n211 );
buf ( n68831 , n68830 );
buf ( n2693 , DFF_rd_reg_Q );
buf ( n2694 , n2693 );
buf ( n2695 , DFF_wr_reg_Q );
buf ( n2696 , n2695 );
buf ( n2697 , n175 );
buf ( n2698 , 1'b0 );
not ( n68838 , n68635 );
not ( n68839 , n68838 );
buf ( n68840 , n68839 );
buf ( n68841 , n68634 );
buf ( n2703 , n63 );
not ( n68843 , n2703 );
not ( n68844 , n68843 );
not ( n68845 , n68844 );
buf ( n68846 , n36 );
not ( n68847 , n68846 );
not ( n68848 , n68847 );
buf ( n2710 , n37 );
not ( n68850 , n2710 );
not ( n68851 , n68850 );
not ( n68852 , n68851 );
not ( n68853 , n68852 );
nor ( n68854 , n68848 , n68853 );
buf ( n68855 , n39 );
not ( n68856 , n68855 );
not ( n68857 , n68856 );
not ( n68858 , n68857 );
not ( n68859 , n68858 );
buf ( n68860 , n38 );
not ( n68861 , n68860 );
not ( n68862 , n68861 );
not ( n68863 , n68862 );
not ( n68864 , n68863 );
nor ( n68865 , n68859 , n68864 );
nand ( n68866 , n68854 , n68865 );
buf ( n2728 , n32 );
not ( n68868 , n2728 );
buf ( n68869 , n33 );
not ( n68870 , n68869 );
nand ( n68871 , n68868 , n68870 );
not ( n68872 , n68871 );
buf ( n2734 , n34 );
not ( n68874 , n2734 );
not ( n68875 , n68874 );
buf ( n68876 , n35 );
not ( n68877 , n68876 );
not ( n68878 , n68877 );
nor ( n68879 , n68875 , n68878 );
nand ( n68880 , n68872 , n68879 );
or ( n68881 , n68866 , n68880 );
not ( n68882 , n68881 );
buf ( n2744 , n41 );
not ( n68884 , n2744 );
buf ( n68885 , n40 );
not ( n68886 , n68885 );
not ( n68887 , n68886 );
not ( n68888 , n68887 );
nand ( n68889 , n68884 , n68888 );
buf ( n68890 , n43 );
not ( n68891 , n68890 );
buf ( n2753 , n42 );
not ( n68893 , n2753 );
nand ( n68894 , n68891 , n68893 );
nor ( n68895 , n68889 , n68894 );
nand ( n68896 , n68882 , n68895 );
buf ( n2758 , n44 );
and ( n68898 , n68896 , n2758 );
not ( n68899 , n68896 );
not ( n68900 , n2758 );
and ( n68901 , n68899 , n68900 );
nor ( n68902 , n68898 , n68901 );
not ( n68903 , n68902 );
not ( n68904 , n68903 );
not ( n68905 , n68904 );
or ( n68906 , n68845 , n68905 );
nand ( n68907 , n68843 , n2758 );
nand ( n68908 , n68906 , n68907 );
not ( n68909 , n68908 );
not ( n68910 , n68909 );
not ( n68911 , n68843 );
not ( n68912 , n68911 );
buf ( n2774 , n47 );
not ( n68914 , n2774 );
not ( n68915 , n68914 );
not ( n68916 , n68880 );
not ( n68917 , n68866 );
nand ( n68918 , n68916 , n68917 );
not ( n68919 , n68918 );
buf ( n68920 , n45 );
not ( n68921 , n68920 );
nand ( n68922 , n68921 , n68900 );
buf ( n2784 , n46 );
nor ( n68924 , n68922 , n2784 );
and ( n68925 , n68895 , n68924 );
nand ( n68926 , n68919 , n68925 );
not ( n68927 , n68926 );
or ( n68928 , n68915 , n68927 );
or ( n68929 , n68926 , n68914 );
nand ( n68930 , n68928 , n68929 );
not ( n68931 , n68930 );
or ( n68932 , n68912 , n68931 );
nand ( n68933 , n68843 , n2774 );
nand ( n68934 , n68932 , n68933 );
nor ( n68935 , n68910 , n68934 );
not ( n68936 , n68844 );
not ( n68937 , n68895 );
nor ( n68938 , n68937 , n2758 );
nand ( n68939 , n68919 , n68938 );
and ( n68940 , n68939 , n68920 );
not ( n68941 , n68939 );
and ( n68942 , n68941 , n68921 );
nor ( n68943 , n68940 , n68942 );
not ( n68944 , n68943 );
or ( n68945 , n68936 , n68944 );
nand ( n68946 , n68843 , n68920 );
nand ( n68947 , n68945 , n68946 );
not ( n68948 , n68947 );
not ( n68949 , n68948 );
not ( n68950 , n68844 );
nor ( n68951 , n68937 , n68922 );
nand ( n68952 , n68919 , n68951 );
and ( n68953 , n68952 , n2784 );
not ( n68954 , n68952 );
not ( n68955 , n2784 );
and ( n68956 , n68954 , n68955 );
nor ( n68957 , n68953 , n68956 );
not ( n68958 , n68957 );
or ( n68959 , n68950 , n68958 );
nand ( n68960 , n68843 , n2784 );
nand ( n68961 , n68959 , n68960 );
nor ( n68962 , n68949 , n68961 );
not ( n68963 , n68844 );
not ( n68964 , n68893 );
nor ( n68965 , n68964 , n68889 );
nand ( n68966 , n68882 , n68965 );
not ( n68967 , n68891 );
and ( n68968 , n68966 , n68967 );
not ( n68969 , n68966 );
and ( n68970 , n68969 , n68891 );
nor ( n68971 , n68968 , n68970 );
not ( n68972 , n68971 );
not ( n68973 , n68972 );
not ( n68974 , n68973 );
or ( n68975 , n68963 , n68974 );
nand ( n68976 , n68843 , n68890 );
nand ( n68977 , n68975 , n68976 );
not ( n68978 , n68977 );
not ( n68979 , n68887 );
not ( n68980 , n68843 );
or ( n68981 , n68979 , n68980 );
not ( n68982 , n68887 );
not ( n68983 , n68882 );
or ( n68984 , n68982 , n68983 );
or ( n68985 , n68919 , n68887 );
nand ( n68986 , n68984 , n68985 );
nand ( n68987 , n68986 , n2703 );
nand ( n68988 , n68981 , n68987 );
and ( n68989 , n68843 , n68857 );
not ( n68990 , n68843 );
not ( n68991 , n68859 );
not ( n68992 , n68991 );
not ( n68993 , n68852 );
nor ( n68994 , n68993 , n68848 );
not ( n68995 , n68994 );
nor ( n68996 , n68995 , n68864 );
not ( n68997 , n68878 );
not ( n68998 , n68869 );
not ( n68999 , n2728 );
not ( n69000 , n68875 );
and ( n69001 , n68997 , n68998 , n68999 , n69000 );
nand ( n69002 , n68996 , n69001 );
not ( n69003 , n69002 );
or ( n69004 , n68992 , n69003 );
nand ( n69005 , n69001 , n68996 );
or ( n69006 , n69005 , n68991 );
nand ( n69007 , n69004 , n69006 );
and ( n69008 , n68990 , n69007 );
nor ( n69009 , n68989 , n69008 );
not ( n69010 , n69009 );
not ( n69011 , n69010 );
and ( n69012 , n68843 , n68851 );
not ( n69013 , n68843 );
not ( n69014 , n68993 );
not ( n69015 , n69014 );
not ( n69016 , n68848 );
nand ( n69017 , n69001 , n69016 );
not ( n69018 , n69017 );
or ( n69019 , n69015 , n69018 );
nand ( n69020 , n69001 , n69016 );
or ( n69021 , n69020 , n69014 );
nand ( n69022 , n69019 , n69021 );
and ( n69023 , n69013 , n69022 );
nor ( n69024 , n69012 , n69023 );
not ( n69025 , n69024 );
not ( n69026 , n69025 );
nand ( n69027 , n69011 , n69026 );
nor ( n69028 , n68988 , n69027 );
and ( n69029 , n68978 , n69028 );
nand ( n69030 , n68935 , n68962 , n69029 );
not ( n69031 , n69030 );
not ( n69032 , n68844 );
not ( n69033 , n68893 );
not ( n69034 , n68889 );
nand ( n69035 , n69034 , n68882 );
not ( n69036 , n69035 );
or ( n69037 , n69033 , n69036 );
or ( n69038 , n69035 , n68893 );
nand ( n69039 , n69037 , n69038 );
not ( n69040 , n69039 );
not ( n69041 , n69040 );
not ( n69042 , n69041 );
or ( n69043 , n69032 , n69042 );
nand ( n69044 , n68843 , n2753 );
nand ( n69045 , n69043 , n69044 );
not ( n69046 , n69045 );
and ( n69047 , n68843 , n68862 );
not ( n69048 , n68843 );
not ( n69049 , n68864 );
not ( n69050 , n69049 );
nand ( n69051 , n69001 , n68994 );
not ( n69052 , n69051 );
or ( n69053 , n69050 , n69052 );
nand ( n69054 , n69001 , n68994 );
or ( n69055 , n69054 , n69049 );
nand ( n69056 , n69053 , n69055 );
and ( n69057 , n69048 , n69056 );
nor ( n69058 , n69047 , n69057 );
not ( n69059 , n69058 );
not ( n69060 , n2703 );
and ( n69061 , n69060 , n68878 );
not ( n69062 , n69060 );
not ( n69063 , n69000 );
nor ( n69064 , n69063 , n68871 );
and ( n69065 , n69064 , n68997 );
not ( n69066 , n69064 );
not ( n69067 , n68997 );
and ( n69068 , n69066 , n69067 );
nor ( n69069 , n69065 , n69068 );
and ( n69070 , n69062 , n69069 );
nor ( n69071 , n69061 , n69070 );
not ( n69072 , n69071 );
not ( n69073 , n69072 );
not ( n69074 , n69016 );
not ( n69075 , n68880 );
or ( n69076 , n69074 , n69075 );
or ( n69077 , n69016 , n68880 );
nand ( n69078 , n69076 , n69077 );
and ( n69079 , n2703 , n69078 );
not ( n69080 , n2703 );
and ( n69081 , n69080 , n68848 );
nor ( n69082 , n69079 , n69081 );
not ( n69083 , n69082 );
not ( n69084 , n69083 );
not ( n69085 , n2703 );
not ( n69086 , n69000 );
not ( n69087 , n68871 );
or ( n69088 , n69086 , n69087 );
or ( n69089 , n68871 , n69000 );
nand ( n69090 , n69088 , n69089 );
not ( n69091 , n69090 );
or ( n69092 , n69085 , n69091 );
not ( n69093 , n2703 );
nand ( n69094 , n69093 , n68875 );
nand ( n69095 , n69092 , n69094 );
not ( n69096 , n2703 );
not ( n69097 , n68998 );
not ( n69098 , n69097 );
not ( n69099 , n68999 );
or ( n69100 , n69098 , n69099 );
or ( n69101 , n69097 , n68999 );
nand ( n69102 , n69100 , n69101 );
not ( n69103 , n69102 );
or ( n69104 , n69096 , n69103 );
nand ( n69105 , n69093 , n68869 );
nand ( n69106 , n69104 , n69105 );
not ( n69107 , n69106 );
not ( n69108 , n2728 );
nand ( n69109 , n69107 , n69108 );
nor ( n69110 , n69095 , n69109 );
nand ( n69111 , n69073 , n69084 , n69110 );
nor ( n69112 , n69059 , n69111 );
and ( n69113 , n69046 , n69112 );
not ( n69114 , n68844 );
nand ( n69115 , n68919 , n68888 );
and ( n69116 , n69115 , n2744 );
not ( n69117 , n69115 );
and ( n69118 , n69117 , n68884 );
nor ( n69119 , n69116 , n69118 );
not ( n69120 , n69119 );
or ( n69121 , n69114 , n69120 );
nand ( n69122 , n68843 , n2744 );
nand ( n69123 , n69121 , n69122 );
not ( n69124 , n69123 );
not ( n69125 , n68844 );
nand ( n69126 , n68893 , n68863 );
nand ( n69127 , n68891 , n68858 );
nor ( n69128 , n69126 , n69127 );
not ( n69129 , n68871 );
nor ( n69130 , n68887 , n68848 );
nand ( n69131 , n69128 , n69129 , n69130 );
nor ( n69132 , n68875 , n2758 );
nor ( n69133 , n68920 , n68878 );
nor ( n69134 , n2774 , n2784 );
nor ( n69135 , n2744 , n68851 );
nand ( n69136 , n69132 , n69133 , n69134 , n69135 );
nor ( n69137 , n69131 , n69136 );
buf ( n69138 , n49 );
buf ( n3000 , n48 );
not ( n69140 , n3000 );
not ( n69141 , n69140 );
nor ( n69142 , n69138 , n69141 );
not ( n69143 , n69142 );
not ( n69144 , n69143 );
nand ( n69145 , n69137 , n69144 );
buf ( n69146 , n50 );
not ( n69147 , n69146 );
not ( n69148 , n69147 );
and ( n69149 , n69145 , n69148 );
not ( n69150 , n69145 );
not ( n69151 , n69148 );
and ( n69152 , n69150 , n69151 );
nor ( n69153 , n69149 , n69152 );
not ( n69154 , n69153 );
or ( n69155 , n69125 , n69154 );
nand ( n69156 , n68843 , n69148 );
nand ( n69157 , n69155 , n69156 );
not ( n69158 , n69157 );
and ( n69159 , n69124 , n69158 );
not ( n69160 , n68844 );
not ( n69161 , n69137 );
nor ( n69162 , n69161 , n69141 );
or ( n69163 , n69162 , n69138 );
nand ( n69164 , n69133 , n69134 , n69130 , n69135 );
not ( n69165 , n69164 );
not ( n69166 , n69128 );
not ( n69167 , n69141 );
nand ( n69168 , n69167 , n68999 , n68998 , n69138 );
not ( n69169 , n69132 );
nor ( n69170 , n69166 , n69168 , n69169 );
nand ( n69171 , n69165 , n69170 );
nand ( n69172 , n69163 , n69171 );
not ( n69173 , n69172 );
or ( n69174 , n69160 , n69173 );
nand ( n69175 , n68843 , n69138 );
nand ( n69176 , n69174 , n69175 );
not ( n69177 , n69176 );
not ( n69178 , n69141 );
not ( n69179 , n68843 );
or ( n69180 , n69178 , n69179 );
not ( n69181 , n69141 );
not ( n69182 , n69137 );
or ( n69183 , n69181 , n69182 );
or ( n69184 , n69137 , n69141 );
nand ( n69185 , n69183 , n69184 );
nand ( n69186 , n69185 , n2703 );
nand ( n69187 , n69180 , n69186 );
not ( n69188 , n69187 );
and ( n69189 , n69177 , n69188 );
nand ( n69190 , n69113 , n69159 , n69189 );
not ( n69191 , n69190 );
and ( n69192 , n69031 , n69191 );
not ( n69193 , n69161 );
buf ( n69194 , n57 );
buf ( n69195 , n56 );
nor ( n69196 , n69194 , n69195 );
buf ( n3058 , n58 );
buf ( n3059 , n59 );
nor ( n69199 , n3058 , n3059 );
nand ( n69200 , n69196 , n69199 );
not ( n69201 , n69200 );
buf ( n69202 , n61 );
buf ( n69203 , n60 );
or ( n69204 , n69202 , n69203 );
buf ( n3066 , n62 );
nor ( n69206 , n69204 , n3066 );
nand ( n69207 , n69201 , n69206 );
buf ( n69208 , n53 );
not ( n69209 , n69208 );
not ( n69210 , n69209 );
buf ( n69211 , n51 );
nor ( n69212 , n69210 , n69211 );
buf ( n69213 , n54 );
nor ( n69214 , n69213 , n69141 );
buf ( n69215 , n55 );
nor ( n69216 , n69215 , n69138 );
buf ( n69217 , n52 );
not ( n69218 , n69217 );
not ( n69219 , n69218 );
nor ( n69220 , n69219 , n69148 );
nand ( n69221 , n69212 , n69214 , n69216 , n69220 );
nor ( n69222 , n69207 , n69221 );
nand ( n69223 , n69193 , n69222 );
and ( n69224 , n69223 , n2703 );
not ( n69225 , n69223 );
not ( n69226 , n2703 );
and ( n69227 , n69225 , n69226 );
nor ( n69228 , n69224 , n69227 );
nand ( n69229 , n69228 , n68844 );
not ( n69230 , n69229 );
not ( n69231 , n69230 );
nor ( n69232 , n69192 , n69231 );
not ( n69233 , n69211 );
not ( n69234 , n68843 );
or ( n69235 , n69233 , n69234 );
nor ( n69236 , n69143 , n69148 );
nand ( n69237 , n69137 , n69236 );
xor ( n69238 , n69237 , n69211 );
nand ( n69239 , n69238 , n68844 );
nand ( n69240 , n69235 , n69239 );
not ( n69241 , n69240 );
not ( n69242 , n68911 );
nor ( n69243 , n69148 , n69211 );
nand ( n69244 , n69142 , n69243 );
not ( n69245 , n69244 );
nand ( n69246 , n69245 , n69137 );
and ( n69247 , n69246 , n69219 );
not ( n69248 , n69246 );
not ( n69249 , n69219 );
and ( n69250 , n69248 , n69249 );
nor ( n69251 , n69247 , n69250 );
not ( n69252 , n69251 );
or ( n69253 , n69242 , n69252 );
not ( n69254 , n68844 );
nand ( n69255 , n69254 , n69219 );
nand ( n69256 , n69253 , n69255 );
not ( n69257 , n69256 );
not ( n69258 , n68911 );
nor ( n69259 , n69244 , n69219 );
nand ( n69260 , n69137 , n69259 );
xor ( n69261 , n69260 , n69210 );
not ( n69262 , n69261 );
or ( n69263 , n69258 , n69262 );
nand ( n69264 , n68843 , n69210 );
nand ( n69265 , n69263 , n69264 );
not ( n69266 , n69265 );
not ( n69267 , n68911 );
nor ( n69268 , n69210 , n69219 );
not ( n69269 , n69268 );
nor ( n69270 , n69269 , n69244 );
nand ( n69271 , n69137 , n69270 );
not ( n69272 , n69213 );
xnor ( n69273 , n69271 , n69272 );
not ( n69274 , n69273 );
or ( n69275 , n69267 , n69274 );
nand ( n69276 , n68843 , n69213 );
nand ( n69277 , n69275 , n69276 );
not ( n69278 , n69277 );
and ( n69279 , n69241 , n69257 , n69266 , n69278 );
not ( n69280 , n68844 );
nand ( n69281 , n69268 , n69272 );
nor ( n69282 , n69244 , n69281 );
nand ( n69283 , n69137 , n69282 );
not ( n69284 , n69215 );
xnor ( n69285 , n69283 , n69284 );
not ( n69286 , n69285 );
or ( n69287 , n69280 , n69286 );
nand ( n69288 , n69254 , n69215 );
nand ( n69289 , n69287 , n69288 );
not ( n69290 , n68911 );
nor ( n69291 , n69221 , n69195 );
nand ( n69292 , n69137 , n69291 );
not ( n69293 , n69194 );
xnor ( n69294 , n69292 , n69293 );
not ( n69295 , n69294 );
or ( n69296 , n69290 , n69295 );
nand ( n69297 , n68843 , n69194 );
nand ( n69298 , n69296 , n69297 );
not ( n69299 , n68911 );
not ( n69300 , n69195 );
not ( n69301 , n69300 );
not ( n69302 , n69221 );
nand ( n69303 , n69302 , n69137 );
not ( n69304 , n69303 );
or ( n69305 , n69301 , n69304 );
or ( n69306 , n69303 , n69300 );
nand ( n69307 , n69305 , n69306 );
not ( n69308 , n69307 );
or ( n69309 , n69299 , n69308 );
nand ( n69310 , n68843 , n69195 );
nand ( n69311 , n69309 , n69310 );
or ( n69312 , n69289 , n69298 , n69311 );
not ( n69313 , n68844 );
not ( n69314 , n69196 );
nor ( n69315 , n69314 , n69221 );
nand ( n69316 , n69137 , n69315 );
not ( n69317 , n3058 );
xnor ( n69318 , n69316 , n69317 );
not ( n69319 , n69318 );
not ( n69320 , n69319 );
not ( n69321 , n69320 );
or ( n69322 , n69313 , n69321 );
nand ( n69323 , n68843 , n3058 );
nand ( n69324 , n69322 , n69323 );
nor ( n69325 , n69312 , n69324 );
and ( n69326 , n69279 , n69325 );
nor ( n69327 , n69326 , n69231 );
nor ( n69328 , n69232 , n69327 );
not ( n69329 , n69328 );
not ( n69330 , n3059 );
not ( n69331 , n69254 );
or ( n69332 , n69330 , n69331 );
nand ( n69333 , n69196 , n69317 );
nor ( n69334 , n69221 , n69333 );
nand ( n69335 , n69137 , n69334 );
xor ( n69336 , n69335 , n3059 );
nand ( n69337 , n69336 , n68844 );
nand ( n69338 , n69332 , n69337 );
nand ( n69339 , n69329 , n69338 );
and ( n69340 , n68843 , n69203 );
not ( n69341 , n68843 );
nor ( n69342 , n69221 , n69200 );
nand ( n69343 , n69137 , n69342 );
not ( n69344 , n69203 );
not ( n69345 , n69344 );
and ( n69346 , n69343 , n69345 );
not ( n69347 , n69343 );
and ( n69348 , n69347 , n69344 );
nor ( n69349 , n69346 , n69348 );
and ( n69350 , n69341 , n69349 );
nor ( n69351 , n69340 , n69350 );
not ( n69352 , n69351 );
not ( n69353 , n69352 );
and ( n69354 , n69339 , n69353 );
not ( n69355 , n69339 );
and ( n69356 , n69355 , n69352 );
nor ( n69357 , n69354 , n69356 );
not ( n69358 , n69357 );
not ( n69359 , n69358 );
nand ( n69360 , n69186 , n69009 );
not ( n69361 , n69360 );
not ( n69362 , n68987 );
nand ( n69363 , n69058 , n69024 );
nor ( n69364 , n69362 , n69363 );
nor ( n69365 , n68930 , n69294 );
nand ( n69366 , n69361 , n69364 , n69365 );
nor ( n69367 , n69285 , n2728 );
nand ( n69368 , n69367 , n69319 , n69040 , n68903 );
nor ( n69369 , n69366 , n69368 );
nor ( n69370 , n69307 , n69261 );
nor ( n69371 , n69251 , n69153 );
nand ( n69372 , n69351 , n69337 , n69370 , n69371 );
not ( n69373 , n69372 );
not ( n69374 , n69119 );
nor ( n69375 , n69095 , n69106 );
and ( n69376 , n69082 , n69071 , n69375 );
nand ( n69377 , n69239 , n69374 , n68972 , n69376 );
nor ( n69378 , n68943 , n68957 );
nor ( n69379 , n69273 , n69172 );
nand ( n69380 , n69378 , n69379 );
nor ( n69381 , n69377 , n69380 );
nand ( n69382 , n69369 , n69373 , n69381 );
nand ( n69383 , n69201 , n69344 );
nor ( n69384 , n69383 , n69221 );
nand ( n69385 , n69193 , n69384 );
xor ( n69386 , n69385 , n69202 );
and ( n69387 , n69386 , n68911 );
and ( n69388 , n68843 , n69202 );
nor ( n69389 , n69387 , n69388 );
nor ( n69390 , n69389 , n69229 );
nand ( n69391 , n69382 , n69390 );
not ( n69392 , n69391 );
not ( n69393 , n69204 );
nand ( n69394 , n69393 , n69201 );
nor ( n69395 , n69394 , n69221 );
nand ( n69396 , n69193 , n69395 );
xor ( n69397 , n69396 , n3066 );
nand ( n69398 , n69397 , n68911 );
nand ( n69399 , n68843 , n3066 );
nand ( n69400 , n69398 , n69399 );
not ( n69401 , n69400 );
and ( n69402 , n69392 , n69401 );
and ( n69403 , n69391 , n69400 );
nor ( n69404 , n69402 , n69403 );
not ( n69405 , n69404 );
nand ( n69406 , n69382 , n69230 );
and ( n69407 , n69406 , n69389 );
not ( n69408 , n69406 );
not ( n69409 , n69389 );
and ( n69410 , n69408 , n69409 );
nor ( n69411 , n69407 , n69410 );
not ( n69412 , n69411 );
nand ( n69413 , n69405 , n69412 );
not ( n69414 , n69413 );
buf ( n3276 , n165 );
nand ( n69416 , n69414 , n3276 );
not ( n69417 , n69404 );
nor ( n69418 , n69412 , n69417 );
not ( n69419 , n69418 );
not ( n69420 , n69419 );
buf ( n3282 , n101 );
nand ( n69422 , n69420 , n3282 );
not ( n69423 , n69411 );
not ( n69424 , n69423 );
nand ( n69425 , n69405 , n69424 );
not ( n69426 , n69425 );
buf ( n3288 , n72 );
nand ( n69428 , n69426 , n3288 );
nand ( n69429 , n69404 , n69423 );
not ( n69430 , n69429 );
buf ( n3292 , n133 );
not ( n69432 , n3292 );
not ( n69433 , n69432 );
nand ( n69434 , n69430 , n69433 );
nand ( n69435 , n69416 , n69422 , n69428 , n69434 );
not ( n69436 , n69413 );
buf ( n69437 , n162 );
nand ( n69438 , n69436 , n69437 );
not ( n69439 , n69419 );
buf ( n3301 , n98 );
nand ( n69441 , n69439 , n3301 );
not ( n69442 , n69425 );
buf ( n3304 , n69 );
nand ( n69444 , n69442 , n3304 );
nand ( n69445 , n69404 , n69412 );
not ( n69446 , n69445 );
buf ( n69447 , n130 );
not ( n69448 , n69447 );
not ( n69449 , n69448 );
nand ( n69450 , n69446 , n69449 );
nand ( n69451 , n69438 , n69441 , n69444 , n69450 );
nand ( n69452 , n69435 , n69451 );
not ( n69453 , n69404 );
nor ( n69454 , n69453 , n69412 );
buf ( n3316 , n102 );
nand ( n69456 , n69454 , n3316 );
nand ( n69457 , n69417 , n69423 );
not ( n69458 , n69457 );
buf ( n3320 , n166 );
nand ( n69460 , n69458 , n3320 );
nand ( n69461 , n69424 , n69453 );
not ( n69462 , n69461 );
buf ( n3324 , n73 );
nand ( n69464 , n69462 , n3324 );
not ( n69465 , n69429 );
buf ( n3327 , n134 );
not ( n69467 , n3327 );
not ( n69468 , n69467 );
nand ( n69469 , n69465 , n69468 );
nand ( n69470 , n69456 , n69460 , n69464 , n69469 );
not ( n69471 , n69461 );
nand ( n69472 , n69470 , n69471 );
nor ( n69473 , n69452 , n69472 );
not ( n69474 , n69445 );
buf ( n3336 , n131 );
not ( n69476 , n3336 );
not ( n69477 , n69476 );
nand ( n69478 , n69474 , n69477 );
not ( n69479 , n69418 );
not ( n69480 , n69479 );
buf ( n3342 , n99 );
nand ( n69482 , n69480 , n3342 );
buf ( n3344 , n70 );
nand ( n69484 , n69426 , n3344 );
buf ( n3346 , n163 );
nand ( n69486 , n69414 , n3346 );
nand ( n69487 , n69478 , n69482 , n69484 , n69486 );
not ( n69488 , n69413 );
buf ( n3350 , n164 );
nand ( n69490 , n69488 , n3350 );
not ( n69491 , n69479 );
buf ( n69492 , n100 );
nand ( n69493 , n69491 , n69492 );
not ( n69494 , n69425 );
buf ( n3356 , n71 );
nand ( n69496 , n69494 , n3356 );
not ( n69497 , n69445 );
buf ( n3359 , n132 );
not ( n69499 , n3359 );
not ( n69500 , n69499 );
nand ( n69501 , n69497 , n69500 );
nand ( n69502 , n69490 , n69493 , n69496 , n69501 );
and ( n69503 , n69487 , n69502 );
nand ( n69504 , n69473 , n69503 );
not ( n69505 , n69504 );
not ( n69506 , n69457 );
buf ( n69507 , n170 );
nand ( n69508 , n69506 , n69507 );
buf ( n69509 , n106 );
nand ( n69510 , n69454 , n69509 );
not ( n69511 , n69461 );
buf ( n69512 , n77 );
nand ( n69513 , n69511 , n69512 );
not ( n69514 , n69429 );
buf ( n69515 , n138 );
not ( n69516 , n69515 );
not ( n69517 , n69516 );
nand ( n69518 , n69514 , n69517 );
nand ( n69519 , n69508 , n69510 , n69513 , n69518 );
buf ( n69520 , n76 );
nand ( n69521 , n69511 , n69520 );
buf ( n69522 , n169 );
nand ( n69523 , n69506 , n69522 );
buf ( n69524 , n105 );
nand ( n69525 , n69454 , n69524 );
not ( n69526 , n69429 );
buf ( n69527 , n137 );
not ( n69528 , n69527 );
not ( n69529 , n69528 );
nand ( n69530 , n69526 , n69529 );
nand ( n69531 , n69521 , n69523 , n69525 , n69530 );
nand ( n69532 , n69519 , n69531 );
buf ( n69533 , n168 );
nand ( n69534 , n69458 , n69533 );
buf ( n69535 , n104 );
nand ( n69536 , n69454 , n69535 );
buf ( n69537 , n75 );
nand ( n69538 , n69462 , n69537 );
buf ( n69539 , n136 );
not ( n69540 , n69539 );
not ( n69541 , n69540 );
nand ( n69542 , n69430 , n69541 );
nand ( n69543 , n69534 , n69536 , n69538 , n69542 );
buf ( n3405 , n167 );
nand ( n69545 , n69458 , n3405 );
buf ( n69546 , n103 );
nand ( n69547 , n69454 , n69546 );
not ( n69548 , n69461 );
buf ( n69549 , n74 );
nand ( n69550 , n69548 , n69549 );
buf ( n3412 , n135 );
nand ( n69552 , n69430 , n3412 );
nand ( n69553 , n69545 , n69547 , n69550 , n69552 );
nand ( n69554 , n69543 , n69553 );
nor ( n69555 , n69532 , n69554 );
not ( n69556 , n69457 );
not ( n69557 , n69556 );
buf ( n69558 , n172 );
not ( n69559 , n69558 );
nor ( n69560 , n69557 , n69559 );
not ( n69561 , n69454 );
buf ( n69562 , n108 );
not ( n69563 , n69562 );
nor ( n69564 , n69561 , n69563 );
nor ( n69565 , n69560 , n69564 );
not ( n69566 , n69461 );
buf ( n69567 , n79 );
and ( n69568 , n69566 , n69567 );
not ( n69569 , n69430 );
buf ( n69570 , n140 );
not ( n69571 , n69570 );
not ( n69572 , n69571 );
not ( n69573 , n69572 );
nor ( n69574 , n69569 , n69573 );
nor ( n69575 , n69568 , n69574 );
nand ( n69576 , n69565 , n69575 );
buf ( n69577 , n171 );
nand ( n69578 , n69506 , n69577 );
buf ( n69579 , n107 );
nand ( n69580 , n69454 , n69579 );
buf ( n3442 , n78 );
nand ( n69582 , n69511 , n3442 );
buf ( n69583 , n139 );
not ( n69584 , n69583 );
not ( n69585 , n69584 );
nand ( n69586 , n69526 , n69585 );
nand ( n69587 , n69578 , n69580 , n69582 , n69586 );
nand ( n69588 , n69576 , n69587 );
buf ( n3450 , n173 );
nand ( n69590 , n69556 , n3450 );
buf ( n69591 , n109 );
nand ( n69592 , n69454 , n69591 );
buf ( n3454 , n80 );
nand ( n69594 , n69426 , n3454 );
buf ( n69595 , n141 );
not ( n69596 , n69595 );
not ( n69597 , n69596 );
nand ( n69598 , n69474 , n69597 );
nand ( n69599 , n69590 , n69592 , n69594 , n69598 );
not ( n69600 , n69599 );
nor ( n69601 , n69588 , n69600 );
nand ( n69602 , n69505 , n69555 , n69601 );
buf ( n69603 , n81 );
nand ( n69604 , n69471 , n69603 );
buf ( n3466 , n174 );
nand ( n69606 , n69414 , n3466 );
buf ( n69607 , n110 );
nand ( n69608 , n69420 , n69607 );
buf ( n3470 , n142 );
not ( n69610 , n3470 );
not ( n69611 , n69610 );
nand ( n69612 , n69474 , n69611 );
nand ( n69613 , n69604 , n69606 , n69608 , n69612 );
not ( n69614 , n69613 );
and ( n69615 , n69602 , n69614 );
not ( n69616 , n69602 );
and ( n69617 , n69616 , n69613 );
nor ( n69618 , n69615 , n69617 );
not ( n69619 , n69618 );
not ( n69620 , n69619 );
and ( n69621 , n69359 , n69620 );
not ( n69622 , n69359 );
nand ( n69623 , n69502 , n69553 , n69487 , n69543 );
nor ( n69624 , n69623 , n69588 );
nand ( n69625 , n69613 , n69599 );
nor ( n69626 , n69532 , n69625 );
and ( n69627 , n69624 , n69626 , n69473 );
buf ( n3489 , n143 );
not ( n69629 , n3489 );
not ( n69630 , n69629 );
nand ( n69631 , n69526 , n69630 );
not ( n69632 , n69458 );
not ( n69633 , n69632 );
nand ( n69634 , n69633 , n2697 );
not ( n69635 , n69454 );
not ( n69636 , n69635 );
buf ( n3498 , n111 );
nand ( n69638 , n69636 , n3498 );
buf ( n69639 , n82 );
nand ( n69640 , n69471 , n69639 );
nand ( n69641 , n69631 , n69634 , n69638 , n69640 );
nand ( n69642 , n69627 , n69641 );
buf ( n69643 , n144 );
not ( n69644 , n69643 );
not ( n69645 , n69644 );
nand ( n69646 , n69526 , n69645 );
not ( n69647 , n69454 );
not ( n69648 , n69647 );
buf ( n3510 , n112 );
nand ( n69650 , n69648 , n3510 );
buf ( n69651 , n176 );
nand ( n69652 , n69633 , n69651 );
buf ( n3514 , n83 );
nand ( n69654 , n69471 , n3514 );
nand ( n69655 , n69646 , n69650 , n69652 , n69654 );
not ( n69656 , n69655 );
and ( n69657 , n69642 , n69656 );
not ( n69658 , n69642 );
and ( n69659 , n69658 , n69655 );
nor ( n69660 , n69657 , n69659 );
not ( n69661 , n69660 );
not ( n69662 , n69561 );
buf ( n69663 , n121 );
not ( n69664 , n69663 );
not ( n69665 , n69664 );
and ( n69666 , n69662 , n69665 );
not ( n69667 , n69506 );
buf ( n3529 , n185 );
not ( n69669 , n3529 );
not ( n69670 , n69669 );
not ( n69671 , n69670 );
nor ( n69672 , n69667 , n69671 );
nor ( n69673 , n69666 , n69672 );
buf ( n69674 , n92 );
not ( n69675 , n69674 );
not ( n69676 , n69675 );
and ( n69677 , n69566 , n69676 );
not ( n69678 , n69430 );
buf ( n69679 , n153 );
not ( n69680 , n69679 );
not ( n69681 , n69680 );
not ( n69682 , n69681 );
nor ( n69683 , n69678 , n69682 );
nor ( n69684 , n69677 , n69683 );
nand ( n69685 , n69673 , n69684 );
buf ( n69686 , n186 );
not ( n69687 , n69686 );
not ( n69688 , n69687 );
not ( n69689 , n69688 );
nor ( n69690 , n69457 , n69689 );
buf ( n3552 , n122 );
not ( n69692 , n3552 );
not ( n69693 , n69692 );
not ( n69694 , n69693 );
nor ( n69695 , n69561 , n69694 );
nor ( n69696 , n69690 , n69695 );
buf ( n69697 , n154 );
not ( n69698 , n69697 );
nor ( n69699 , n69569 , n69698 );
buf ( n3561 , n93 );
not ( n69701 , n3561 );
not ( n69702 , n69701 );
not ( n69703 , n69702 );
nor ( n69704 , n69461 , n69703 );
nor ( n69705 , n69699 , n69704 );
nand ( n69706 , n69696 , n69705 );
nand ( n69707 , n69685 , n69706 );
buf ( n3569 , n187 );
not ( n69709 , n3569 );
not ( n69710 , n69709 );
not ( n69711 , n69710 );
nor ( n69712 , n69457 , n69711 );
buf ( n69713 , n123 );
not ( n69714 , n69713 );
not ( n69715 , n69714 );
not ( n69716 , n69715 );
nor ( n69717 , n69561 , n69716 );
nor ( n69718 , n69712 , n69717 );
buf ( n3580 , n94 );
not ( n69720 , n3580 );
not ( n69721 , n69720 );
and ( n69722 , n69566 , n69721 );
buf ( n3584 , n155 );
not ( n69724 , n3584 );
not ( n69725 , n69724 );
not ( n69726 , n69725 );
nor ( n69727 , n69678 , n69726 );
nor ( n69728 , n69722 , n69727 );
nand ( n69729 , n69718 , n69728 );
buf ( n3591 , n156 );
not ( n69731 , n3591 );
not ( n69732 , n69731 );
nand ( n69733 , n69526 , n69732 );
not ( n69734 , n69561 );
buf ( n69735 , n124 );
not ( n69736 , n69735 );
not ( n69737 , n69736 );
nand ( n69738 , n69734 , n69737 );
buf ( n69739 , n188 );
not ( n69740 , n69739 );
not ( n69741 , n69740 );
nand ( n69742 , n69506 , n69741 );
nand ( n69743 , n69733 , n69738 , n69742 );
nand ( n69744 , n69729 , n69743 );
nor ( n69745 , n69707 , n69744 );
not ( n69746 , n69557 );
buf ( n69747 , n182 );
not ( n69748 , n69747 );
not ( n69749 , n69748 );
not ( n69750 , n69749 );
not ( n69751 , n69750 );
and ( n69752 , n69746 , n69751 );
buf ( n69753 , n118 );
not ( n69754 , n69753 );
not ( n69755 , n69754 );
and ( n69756 , n69636 , n69755 );
nor ( n69757 , n69752 , n69756 );
not ( n69758 , n69429 );
buf ( n3620 , n150 );
not ( n69760 , n3620 );
not ( n69761 , n69760 );
not ( n69762 , n69761 );
not ( n69763 , n69762 );
and ( n69764 , n69758 , n69763 );
not ( n69765 , n69461 );
buf ( n69766 , n89 );
and ( n69767 , n69765 , n69766 );
nor ( n69768 , n69764 , n69767 );
nand ( n69769 , n69757 , n69768 );
buf ( n69770 , n88 );
not ( n69771 , n69770 );
not ( n69772 , n69771 );
not ( n69773 , n69772 );
nor ( n69774 , n69461 , n69773 );
buf ( n3636 , n117 );
not ( n69776 , n3636 );
not ( n69777 , n69776 );
not ( n69778 , n69777 );
nor ( n69779 , n69647 , n69778 );
nor ( n69780 , n69774 , n69779 );
buf ( n69781 , n181 );
not ( n69782 , n69781 );
not ( n69783 , n69782 );
not ( n69784 , n69783 );
nor ( n69785 , n69457 , n69784 );
buf ( n69786 , n149 );
not ( n69787 , n69786 );
not ( n69788 , n69787 );
not ( n69789 , n69788 );
nor ( n69790 , n69429 , n69789 );
nor ( n69791 , n69785 , n69790 );
nand ( n69792 , n69780 , n69791 );
nand ( n69793 , n69769 , n69792 );
buf ( n69794 , n146 );
not ( n69795 , n69794 );
not ( n69796 , n69795 );
nand ( n69797 , n69430 , n69796 );
buf ( n69798 , n178 );
nand ( n69799 , n69556 , n69798 );
buf ( n69800 , n114 );
nand ( n69801 , n69636 , n69800 );
buf ( n69802 , n85 );
nand ( n69803 , n69566 , n69802 );
nand ( n69804 , n69797 , n69799 , n69801 , n69803 );
not ( n69805 , n69632 );
buf ( n69806 , n177 );
not ( n69807 , n69806 );
not ( n69808 , n69807 );
and ( n69809 , n69805 , n69808 );
buf ( n69810 , n113 );
and ( n69811 , n69648 , n69810 );
nor ( n69812 , n69809 , n69811 );
buf ( n69813 , n145 );
not ( n69814 , n69813 );
not ( n69815 , n69814 );
not ( n69816 , n69815 );
nor ( n69817 , n69429 , n69816 );
buf ( n69818 , n84 );
not ( n69819 , n69818 );
nor ( n69820 , n69461 , n69819 );
nor ( n69821 , n69817 , n69820 );
nand ( n69822 , n69812 , n69821 );
nand ( n69823 , n69804 , n69822 );
nor ( n69824 , n69793 , n69823 );
nand ( n69825 , n69745 , n69824 );
nand ( n69826 , n69655 , n69641 );
not ( n69827 , n69826 );
not ( n69828 , n69457 );
buf ( n69829 , n184 );
not ( n69830 , n69829 );
not ( n69831 , n69830 );
not ( n69832 , n69831 );
not ( n69833 , n69832 );
and ( n69834 , n69828 , n69833 );
buf ( n69835 , n120 );
not ( n69836 , n69835 );
not ( n69837 , n69836 );
and ( n69838 , n69662 , n69837 );
nor ( n69839 , n69834 , n69838 );
buf ( n69840 , n152 );
not ( n69841 , n69840 );
not ( n69842 , n69841 );
not ( n69843 , n69842 );
nor ( n69844 , n69569 , n69843 );
not ( n69845 , n69566 );
buf ( n3707 , n91 );
not ( n69847 , n3707 );
nor ( n69848 , n69845 , n69847 );
nor ( n69849 , n69844 , n69848 );
nand ( n69850 , n69839 , n69849 );
buf ( n69851 , n86 );
not ( n69852 , n69851 );
nor ( n69853 , n69461 , n69852 );
buf ( n69854 , n115 );
not ( n69855 , n69854 );
not ( n69856 , n69855 );
not ( n69857 , n69856 );
nor ( n69858 , n69635 , n69857 );
nor ( n69859 , n69853 , n69858 );
buf ( n3721 , n179 );
not ( n69861 , n3721 );
not ( n69862 , n69861 );
not ( n69863 , n69862 );
nor ( n69864 , n69457 , n69863 );
buf ( n69865 , n147 );
not ( n69866 , n69865 );
not ( n69867 , n69866 );
not ( n69868 , n69867 );
nor ( n69869 , n69429 , n69868 );
nor ( n69870 , n69864 , n69869 );
nand ( n69871 , n69859 , n69870 );
and ( n69872 , n69850 , n69871 );
not ( n69873 , n69457 );
buf ( n69874 , n180 );
not ( n69875 , n69874 );
not ( n69876 , n69875 );
not ( n69877 , n69876 );
not ( n69878 , n69877 );
and ( n69879 , n69873 , n69878 );
buf ( n69880 , n116 );
not ( n69881 , n69880 );
not ( n69882 , n69881 );
and ( n69883 , n69636 , n69882 );
nor ( n69884 , n69879 , n69883 );
buf ( n69885 , n87 );
not ( n69886 , n69885 );
not ( n69887 , n69886 );
not ( n69888 , n69887 );
nor ( n69889 , n69461 , n69888 );
buf ( n69890 , n148 );
not ( n69891 , n69890 );
not ( n69892 , n69891 );
not ( n69893 , n69892 );
nor ( n69894 , n69429 , n69893 );
nor ( n69895 , n69889 , n69894 );
nand ( n69896 , n69884 , n69895 );
buf ( n69897 , n125 );
not ( n69898 , n69897 );
not ( n69899 , n69898 );
nand ( n69900 , n69662 , n69899 );
not ( n69901 , n69457 );
buf ( n69902 , n189 );
nand ( n69903 , n69901 , n69902 );
buf ( n69904 , n157 );
not ( n69905 , n69904 );
not ( n69906 , n69905 );
nand ( n69907 , n69526 , n69906 );
nand ( n69908 , n69900 , n69903 , n69907 );
and ( n69909 , n69896 , n69908 );
buf ( n3771 , n119 );
not ( n69911 , n3771 );
not ( n69912 , n69911 );
and ( n69913 , n69734 , n69912 );
buf ( n69914 , n183 );
not ( n69915 , n69914 );
not ( n69916 , n69915 );
not ( n69917 , n69916 );
nor ( n69918 , n69667 , n69917 );
nor ( n69919 , n69913 , n69918 );
not ( n69920 , n69526 );
buf ( n69921 , n151 );
not ( n69922 , n69921 );
not ( n69923 , n69922 );
not ( n69924 , n69923 );
nor ( n69925 , n69920 , n69924 );
buf ( n69926 , n90 );
not ( n69927 , n69926 );
not ( n69928 , n69927 );
not ( n69929 , n69928 );
nor ( n69930 , n69461 , n69929 );
nor ( n69931 , n69925 , n69930 );
nand ( n69932 , n69919 , n69931 );
nand ( n69933 , n69827 , n69872 , n69909 , n69932 );
nor ( n69934 , n69825 , n69933 );
nand ( n69935 , n69627 , n69934 );
buf ( n69936 , n126 );
nand ( n69937 , n69734 , n69936 );
buf ( n3799 , n158 );
nand ( n69939 , n69526 , n3799 );
buf ( n69940 , n190 );
nand ( n69941 , n69506 , n69940 );
nand ( n69942 , n69937 , n69939 , n69941 );
not ( n69943 , n69942 );
and ( n69944 , n69935 , n69943 );
not ( n69945 , n69935 );
and ( n69946 , n69945 , n69942 );
nor ( n69947 , n69944 , n69946 );
buf ( n69948 , n66 );
not ( n69949 , n69948 );
not ( n69950 , n69949 );
not ( n69951 , n69950 );
not ( n69952 , n69471 );
or ( n69953 , n69951 , n69952 );
buf ( n3815 , n159 );
nand ( n69955 , n69901 , n3815 );
nand ( n69956 , n69953 , n69955 );
buf ( n69957 , n95 );
not ( n69958 , n69957 );
not ( n69959 , n69636 );
or ( n69960 , n69958 , n69959 );
buf ( n69961 , n127 );
not ( n69962 , n69961 );
not ( n69963 , n69962 );
nand ( n69964 , n69430 , n69963 );
nand ( n69965 , n69960 , n69964 );
nor ( n69966 , n69956 , n69965 );
not ( n69967 , n69966 );
nand ( n69968 , n69947 , n69967 );
not ( n69969 , n69968 );
not ( n69970 , n69969 );
not ( n69971 , n69970 );
not ( n69972 , n69641 );
not ( n69973 , n69627 );
not ( n69974 , n69973 );
or ( n69975 , n69972 , n69974 );
or ( n69976 , n69973 , n69641 );
nand ( n69977 , n69975 , n69976 );
not ( n69978 , n69977 );
not ( n69979 , n69588 );
nand ( n69980 , n69979 , n69505 , n69555 );
xor ( n69981 , n69980 , n69600 );
nand ( n69982 , n69618 , n69981 );
nor ( n69983 , n69978 , n69982 );
not ( n69984 , n69983 );
nand ( n69985 , n69505 , n69555 );
not ( n69986 , n69587 );
and ( n69987 , n69985 , n69986 );
not ( n69988 , n69985 );
and ( n69989 , n69988 , n69587 );
nor ( n69990 , n69987 , n69989 );
not ( n69991 , n69554 );
not ( n69992 , n69991 );
not ( n69993 , n69531 );
nor ( n69994 , n69992 , n69993 );
nand ( n69995 , n69505 , n69994 );
not ( n69996 , n69519 );
and ( n69997 , n69995 , n69996 );
not ( n69998 , n69995 );
and ( n69999 , n69998 , n69519 );
nor ( n70000 , n69997 , n69999 );
nand ( n70001 , n69990 , n70000 );
nand ( n70002 , n69505 , n69553 );
not ( n70003 , n69543 );
and ( n70004 , n70002 , n70003 );
not ( n70005 , n70002 );
and ( n70006 , n70005 , n69543 );
nor ( n70007 , n70004 , n70006 );
nand ( n70008 , n69505 , n69991 );
not ( n70009 , n69531 );
and ( n70010 , n70008 , n70009 );
not ( n70011 , n70008 );
and ( n70012 , n70011 , n69531 );
nor ( n70013 , n70010 , n70012 );
and ( n70014 , n70007 , n70013 );
not ( n70015 , n70014 );
nor ( n70016 , n70001 , n70015 );
nand ( n70017 , n69451 , n69471 );
not ( n70018 , n69487 );
or ( n70019 , n70017 , n70018 );
not ( n70020 , n69502 );
and ( n70021 , n70019 , n70020 );
not ( n70022 , n70019 );
and ( n70023 , n70022 , n69502 );
nor ( n70024 , n70021 , n70023 );
not ( n70025 , n69503 );
or ( n70026 , n70017 , n70025 );
not ( n70027 , n69435 );
and ( n70028 , n70026 , n70027 );
not ( n70029 , n70026 );
and ( n70030 , n70029 , n69435 );
nor ( n70031 , n70028 , n70030 );
nand ( n70032 , n70024 , n70031 );
not ( n70033 , n69487 );
nand ( n70034 , n69451 , n69471 );
not ( n70035 , n70034 );
or ( n70036 , n70033 , n70035 );
or ( n70037 , n70034 , n69487 );
nand ( n70038 , n70036 , n70037 );
or ( n70039 , n69451 , n69471 );
and ( n70040 , n70034 , n70039 );
buf ( n70041 , n67 );
nand ( n70042 , n69471 , n70041 );
buf ( n70043 , n128 );
not ( n70044 , n70043 );
not ( n70045 , n70044 );
nand ( n70046 , n69430 , n70045 );
buf ( n70047 , n96 );
not ( n70048 , n70047 );
not ( n70049 , n70048 );
nand ( n70050 , n69636 , n70049 );
buf ( n70051 , n160 );
nand ( n70052 , n69901 , n70051 );
nand ( n70053 , n70042 , n70046 , n70050 , n70052 );
buf ( n3915 , n68 );
not ( n70055 , n3915 );
not ( n70056 , n69471 );
or ( n70057 , n70055 , n70056 );
buf ( n70058 , n161 );
nand ( n70059 , n69901 , n70058 );
nand ( n70060 , n70057 , n70059 );
buf ( n70061 , n129 );
not ( n70062 , n70061 );
not ( n70063 , n70062 );
not ( n70064 , n70063 );
not ( n70065 , n69430 );
or ( n70066 , n70064 , n70065 );
buf ( n70067 , n97 );
not ( n70068 , n70067 );
not ( n70069 , n70068 );
nand ( n70070 , n69636 , n70069 );
nand ( n70071 , n70066 , n70070 );
nor ( n70072 , n70060 , n70071 );
not ( n70073 , n70072 );
and ( n70074 , n70053 , n70073 );
nand ( n70075 , n70038 , n70040 , n70074 );
nor ( n70076 , n70032 , n70075 );
not ( n70077 , n69553 );
not ( n70078 , n69505 );
not ( n70079 , n70078 );
or ( n70080 , n70077 , n70079 );
or ( n70081 , n70078 , n69553 );
nand ( n70082 , n70080 , n70081 );
not ( n70083 , n69470 );
not ( n70084 , n70034 );
nor ( n70085 , n70025 , n70027 );
nand ( n70086 , n70084 , n70085 );
not ( n70087 , n70086 );
or ( n70088 , n70083 , n70087 );
or ( n70089 , n70086 , n69470 );
nand ( n70090 , n70088 , n70089 );
nand ( n70091 , n70076 , n70082 , n70090 );
not ( n70092 , n70091 );
nand ( n70093 , n69505 , n69555 , n69587 );
not ( n70094 , n69576 );
and ( n70095 , n70093 , n70094 );
not ( n70096 , n70093 );
and ( n70097 , n70096 , n69576 );
nor ( n70098 , n70095 , n70097 );
nand ( n70099 , n70016 , n70092 , n70098 );
not ( n70100 , n70099 );
not ( n70101 , n70100 );
nor ( n70102 , n69984 , n70101 );
nand ( n70103 , n69971 , n70102 );
not ( n70104 , n70103 );
or ( n70105 , n69661 , n70104 );
or ( n70106 , n70103 , n69660 );
nand ( n70107 , n70105 , n70106 );
and ( n70108 , n69622 , n70107 );
nor ( n70109 , n69621 , n70108 );
not ( n70110 , n69298 );
not ( n70111 , n69289 );
not ( n70112 , n69230 );
or ( n70113 , n70111 , n70112 );
not ( n70114 , n69030 );
not ( n70115 , n69190 );
and ( n70116 , n70114 , n70115 );
nor ( n70117 , n70116 , n69231 );
nor ( n70118 , n69279 , n69231 );
nor ( n70119 , n70117 , n70118 );
nand ( n70120 , n70113 , n70119 );
nand ( n70121 , n70120 , n69311 );
nor ( n70122 , n70110 , n70121 );
xor ( n70123 , n70122 , n69324 );
not ( n70124 , n70121 );
not ( n70125 , n69298 );
and ( n70126 , n70124 , n70125 );
and ( n70127 , n70121 , n69298 );
nor ( n70128 , n70126 , n70127 );
and ( n70129 , n70120 , n69311 );
not ( n70130 , n70120 );
not ( n70131 , n69311 );
and ( n70132 , n70130 , n70131 );
nor ( n70133 , n70129 , n70132 );
not ( n70134 , n70133 );
nor ( n70135 , n70128 , n70134 );
nand ( n70136 , n70123 , n70135 );
buf ( n70137 , DFF_state_reg_Q );
not ( n70138 , n70137 );
not ( n70139 , n70138 );
and ( n70140 , n70136 , n70139 );
not ( n70141 , n70140 );
not ( n70142 , n70119 );
not ( n70143 , n69289 );
and ( n70144 , n70142 , n70143 );
and ( n70145 , n70119 , n69289 );
nor ( n70146 , n70144 , n70145 );
not ( n70147 , n70146 );
nor ( n70148 , n70141 , n70147 );
not ( n70149 , n70128 );
not ( n70150 , n70149 );
buf ( n70151 , DFF_B_reg_Q );
not ( n70152 , n70151 );
nand ( n70153 , n70150 , n70152 );
not ( n70154 , n70153 );
not ( n70155 , n70123 );
or ( n70156 , n70154 , n70155 );
nand ( n70157 , n70156 , n70133 );
not ( n70158 , n70133 );
nand ( n70159 , n70158 , n70151 );
nor ( n70160 , n70149 , n70159 );
buf ( n70161 , n64 );
or ( n70162 , n70160 , n70161 );
nand ( n70163 , n70162 , n70123 );
nand ( n70164 , n70157 , n70163 );
not ( n70165 , n70149 );
not ( n70166 , n70123 );
not ( n70167 , n70166 );
or ( n70168 , n70165 , n70167 );
buf ( n70169 , n65 );
not ( n70170 , n70169 );
not ( n70171 , n70170 );
nand ( n70172 , n70133 , n70152 );
not ( n70173 , n70172 );
not ( n70174 , n70159 );
or ( n70175 , n70173 , n70174 );
nand ( n70176 , n70175 , n70150 );
not ( n70177 , n70176 );
or ( n70178 , n70171 , n70177 );
nand ( n70179 , n70178 , n70123 );
nand ( n70180 , n70168 , n70179 );
not ( n70181 , n70180 );
nor ( n70182 , n70164 , n70181 );
nand ( n70183 , n70148 , n70182 );
not ( n70184 , n69241 );
nand ( n70185 , n70117 , n70184 );
nor ( n70186 , n70185 , n69257 );
nand ( n70187 , n70186 , n69265 );
xor ( n70188 , n70187 , n69278 );
not ( n70189 , n69265 );
nor ( n70190 , n70189 , n70186 );
not ( n70191 , n70190 );
not ( n70192 , n69265 );
nand ( n70193 , n70192 , n70186 );
nand ( n70194 , n70191 , n70193 );
nand ( n70195 , n70188 , n70194 );
not ( n70196 , n70195 );
not ( n70197 , n69257 );
not ( n70198 , n70197 );
not ( n70199 , n70185 );
or ( n70200 , n70198 , n70199 );
or ( n70201 , n70185 , n70197 );
nand ( n70202 , n70200 , n70201 );
and ( n70203 , n70117 , n70184 );
not ( n70204 , n70117 );
and ( n70205 , n70204 , n69241 );
nor ( n70206 , n70203 , n70205 );
nor ( n70207 , n70202 , n70206 );
nand ( n70208 , n70196 , n70207 );
nor ( n70209 , n70183 , n70208 );
not ( n70210 , n70209 );
or ( n70211 , n70109 , n70210 );
not ( n70212 , n69641 );
not ( n70213 , n69328 );
not ( n70214 , n69338 );
and ( n70215 , n70213 , n70214 );
and ( n70216 , n69328 , n69338 );
nor ( n70217 , n70215 , n70216 );
and ( n70218 , n69338 , n69353 );
not ( n70219 , n69338 );
and ( n70220 , n70219 , n69352 );
nor ( n70221 , n70218 , n70220 );
nand ( n70222 , n70217 , n70221 );
or ( n70223 , n70222 , n69188 );
nand ( n70224 , n70222 , n68651 );
nand ( n70225 , n70223 , n70224 );
not ( n70226 , n70225 );
or ( n70227 , n70212 , n70226 );
not ( n70228 , n69641 );
not ( n70229 , n70225 );
nand ( n70230 , n70228 , n70229 );
nand ( n70231 , n70227 , n70230 );
not ( n70232 , n70222 );
not ( n70233 , n68934 );
not ( n70234 , n70233 );
and ( n70235 , n70232 , n70234 );
and ( n70236 , n70222 , n2513 );
nor ( n70237 , n70235 , n70236 );
not ( n70238 , n70237 );
not ( n70239 , n70238 );
and ( n70240 , n70239 , n69613 );
nor ( n70241 , n70231 , n70240 );
not ( n70242 , n70241 );
nand ( n70243 , n70231 , n70240 );
nand ( n70244 , n70242 , n70243 );
not ( n70245 , n70244 );
not ( n70246 , n69531 );
not ( n70247 , n70222 );
not ( n70248 , n69045 );
not ( n70249 , n70248 );
and ( n70250 , n70247 , n70249 );
and ( n70251 , n70222 , n2518 );
nor ( n70252 , n70250 , n70251 );
not ( n70253 , n70252 );
not ( n70254 , n70253 );
or ( n70255 , n70246 , n70254 );
not ( n70256 , n70253 );
not ( n70257 , n69531 );
nand ( n70258 , n70256 , n70257 );
nand ( n70259 , n70255 , n70258 );
nor ( n70260 , n70222 , n69124 );
not ( n70261 , n70260 );
nand ( n70262 , n70222 , n2519 );
nand ( n70263 , n70261 , n70262 );
not ( n70264 , n70263 );
and ( n70265 , n69543 , n70264 );
and ( n70266 , n70259 , n70265 );
not ( n70267 , n70266 );
not ( n70268 , n70222 );
not ( n70269 , n68978 );
and ( n70270 , n70268 , n70269 );
and ( n70271 , n70222 , n2517 );
nor ( n70272 , n70270 , n70271 );
not ( n70273 , n70272 );
not ( n70274 , n70273 );
not ( n70275 , n69519 );
or ( n70276 , n70274 , n70275 );
not ( n70277 , n70273 );
not ( n70278 , n69519 );
nand ( n70279 , n70277 , n70278 );
nand ( n70280 , n70276 , n70279 );
nor ( n70281 , n70253 , n70257 );
nor ( n70282 , n70280 , n70281 );
not ( n70283 , n70282 );
not ( n70284 , n70283 );
or ( n70285 , n70267 , n70284 );
nand ( n70286 , n70280 , n70281 );
nand ( n70287 , n70285 , n70286 );
not ( n70288 , n70287 );
not ( n70289 , n69576 );
not ( n70290 , n70289 );
not ( n70291 , n70222 );
not ( n70292 , n68948 );
and ( n70293 , n70291 , n70292 );
and ( n70294 , n70222 , n2515 );
nor ( n70295 , n70293 , n70294 );
not ( n70296 , n70295 );
not ( n70297 , n70296 );
not ( n70298 , n70297 );
or ( n70299 , n70290 , n70298 );
nand ( n70300 , n69576 , n70296 );
nand ( n70301 , n70299 , n70300 );
not ( n70302 , n69587 );
not ( n70303 , n70222 );
not ( n70304 , n68909 );
and ( n70305 , n70303 , n70304 );
and ( n70306 , n70222 , n2516 );
nor ( n70307 , n70305 , n70306 );
not ( n70308 , n70307 );
nor ( n70309 , n70302 , n70308 );
nor ( n70310 , n70301 , n70309 );
not ( n70311 , n69587 );
not ( n70312 , n70308 );
or ( n70313 , n70311 , n70312 );
not ( n70314 , n70308 );
not ( n70315 , n69587 );
nand ( n70316 , n70314 , n70315 );
nand ( n70317 , n70313 , n70316 );
nand ( n70318 , n69519 , n70277 );
not ( n70319 , n70318 );
nor ( n70320 , n70317 , n70319 );
nor ( n70321 , n70310 , n70320 );
not ( n70322 , n69599 );
not ( n70323 , n68961 );
nor ( n70324 , n70222 , n70323 );
not ( n70325 , n70324 );
nand ( n70326 , n70222 , n2514 );
nand ( n70327 , n70325 , n70326 );
not ( n70328 , n70327 );
or ( n70329 , n70322 , n70328 );
not ( n70330 , n69599 );
not ( n70331 , n70327 );
nand ( n70332 , n70330 , n70331 );
nand ( n70333 , n70329 , n70332 );
not ( n70334 , n69576 );
nor ( n70335 , n70334 , n70296 );
nor ( n70336 , n70333 , n70335 );
not ( n70337 , n69613 );
not ( n70338 , n70238 );
or ( n70339 , n70337 , n70338 );
not ( n70340 , n69613 );
nand ( n70341 , n70340 , n70239 );
nand ( n70342 , n70339 , n70341 );
nand ( n70343 , n70331 , n69599 );
not ( n70344 , n70343 );
nor ( n70345 , n70342 , n70344 );
nor ( n70346 , n70336 , n70345 );
and ( n70347 , n70321 , n70346 );
not ( n70348 , n70347 );
or ( n70349 , n70288 , n70348 );
not ( n70350 , n70346 );
nand ( n70351 , n70317 , n70319 );
not ( n70352 , n70351 );
not ( n70353 , n70352 );
not ( n70354 , n70310 );
not ( n70355 , n70354 );
or ( n70356 , n70353 , n70355 );
nand ( n70357 , n70301 , n70309 );
nand ( n70358 , n70356 , n70357 );
not ( n70359 , n70358 );
or ( n70360 , n70350 , n70359 );
not ( n70361 , n70345 );
nand ( n70362 , n70333 , n70335 );
not ( n70363 , n70362 );
and ( n70364 , n70361 , n70363 );
nand ( n70365 , n70342 , n70344 );
not ( n70366 , n70365 );
nor ( n70367 , n70364 , n70366 );
nand ( n70368 , n70360 , n70367 );
not ( n70369 , n70368 );
nand ( n70370 , n70349 , n70369 );
not ( n70371 , n70370 );
nor ( n70372 , n70259 , n70265 );
nor ( n70373 , n70372 , n70282 );
not ( n70374 , n69553 );
not ( n70375 , n68988 );
or ( n70376 , n70222 , n70375 );
nand ( n70377 , n70222 , n68659 );
nand ( n70378 , n70376 , n70377 );
not ( n70379 , n70378 );
or ( n70380 , n70374 , n70379 );
not ( n70381 , n70378 );
not ( n70382 , n69553 );
nand ( n70383 , n70381 , n70382 );
nand ( n70384 , n70380 , n70383 );
not ( n70385 , n70384 );
or ( n70386 , n70222 , n69011 );
nand ( n70387 , n70222 , n68660 );
nand ( n70388 , n70386 , n70387 );
not ( n70389 , n69470 );
nor ( n70390 , n70388 , n70389 );
not ( n70391 , n70390 );
nand ( n70392 , n70385 , n70391 );
xor ( n70393 , n69543 , n70264 );
not ( n70394 , n70393 );
nor ( n70395 , n70378 , n70382 );
not ( n70396 , n70395 );
nand ( n70397 , n70394 , n70396 );
and ( n70398 , n70392 , n70397 );
not ( n70399 , n69487 );
not ( n70400 , n70222 );
not ( n70401 , n69084 );
and ( n70402 , n70400 , n70401 );
and ( n70403 , n70222 , n2524 );
nor ( n70404 , n70402 , n70403 );
not ( n70405 , n70404 );
not ( n70406 , n70405 );
or ( n70407 , n70399 , n70406 );
or ( n70408 , n70405 , n69487 );
nand ( n70409 , n70407 , n70408 );
not ( n70410 , n69471 );
not ( n70411 , n70410 );
not ( n70412 , n69451 );
not ( n70413 , n70412 );
or ( n70414 , n70411 , n70413 );
not ( n70415 , n69072 );
not ( n70416 , n70222 );
not ( n70417 , n70416 );
or ( n70418 , n70415 , n70417 );
nand ( n70419 , n70222 , n68664 );
nand ( n70420 , n70418 , n70419 );
not ( n70421 , n70420 );
nand ( n70422 , n70414 , n70421 );
not ( n70423 , n70412 );
nand ( n70424 , n70423 , n69471 );
nand ( n70425 , n70422 , n70424 );
nor ( n70426 , n70409 , n70425 );
not ( n70427 , n69502 );
not ( n70428 , n69025 );
not ( n70429 , n70416 );
or ( n70430 , n70428 , n70429 );
nand ( n70431 , n70222 , n2523 );
nand ( n70432 , n70430 , n70431 );
not ( n70433 , n70432 );
or ( n70434 , n70427 , n70433 );
not ( n70435 , n70432 );
not ( n70436 , n69502 );
nand ( n70437 , n70435 , n70436 );
nand ( n70438 , n70434 , n70437 );
not ( n70439 , n69487 );
nor ( n70440 , n70439 , n70405 );
nor ( n70441 , n70438 , n70440 );
nor ( n70442 , n70426 , n70441 );
not ( n70443 , n69471 );
not ( n70444 , n69451 );
not ( n70445 , n70444 );
or ( n70446 , n70443 , n70445 );
nand ( n70447 , n69451 , n70410 );
nand ( n70448 , n70446 , n70447 );
and ( n70449 , n70448 , n70421 );
not ( n70450 , n70448 );
and ( n70451 , n70450 , n70420 );
nor ( n70452 , n70449 , n70451 );
not ( n70453 , n70222 );
not ( n70454 , n69095 );
not ( n70455 , n70454 );
and ( n70456 , n70453 , n70455 );
and ( n70457 , n70222 , n68665 );
nor ( n70458 , n70456 , n70457 );
not ( n70459 , n70458 );
not ( n70460 , n70459 );
and ( n70461 , n70073 , n70460 );
nor ( n70462 , n70452 , n70461 );
not ( n70463 , n70462 );
and ( n70464 , n70373 , n70398 , n70442 , n70463 );
not ( n70465 , n70389 );
not ( n70466 , n70388 );
not ( n70467 , n70466 );
or ( n70468 , n70465 , n70467 );
nand ( n70469 , n70388 , n69470 );
nand ( n70470 , n70468 , n70469 );
not ( n70471 , n70222 );
not ( n70472 , n69059 );
not ( n70473 , n70472 );
and ( n70474 , n70471 , n70473 );
and ( n70475 , n70222 , n68661 );
nor ( n70476 , n70474 , n70475 );
not ( n70477 , n70476 );
not ( n70478 , n69435 );
nor ( n70479 , n70477 , n70478 );
nor ( n70480 , n70470 , n70479 );
not ( n70481 , n69435 );
not ( n70482 , n70477 );
or ( n70483 , n70481 , n70482 );
not ( n70484 , n70477 );
nand ( n70485 , n70484 , n70478 );
nand ( n70486 , n70483 , n70485 );
nor ( n70487 , n70432 , n70436 );
nand ( n70488 , n70486 , n70487 );
nor ( n70489 , n70480 , n70488 );
and ( n70490 , n70470 , n70479 );
nor ( n70491 , n70489 , n70490 );
or ( n70492 , n70470 , n70479 );
not ( n70493 , n70486 );
not ( n70494 , n70487 );
nand ( n70495 , n70493 , n70494 );
nand ( n70496 , n70492 , n70495 );
nand ( n70497 , n70491 , n70496 );
not ( n70498 , n70222 );
not ( n70499 , n69107 );
and ( n70500 , n70498 , n70499 );
and ( n70501 , n70222 , n68666 );
nor ( n70502 , n70500 , n70501 );
not ( n70503 , n70502 );
or ( n70504 , n70503 , n70053 );
nand ( n70505 , n70053 , n70503 );
nand ( n70506 , n70504 , n70505 );
nor ( n70507 , n70506 , n69967 );
not ( n70508 , n70460 );
not ( n70509 , n70073 );
not ( n70510 , n70509 );
or ( n70511 , n70508 , n70510 );
nand ( n70512 , n70073 , n70459 );
nand ( n70513 , n70511 , n70512 );
not ( n70514 , n70053 );
nor ( n70515 , n70514 , n70503 );
nor ( n70516 , n70513 , n70515 );
nor ( n70517 , n70507 , n70516 );
nand ( n70518 , n70506 , n69967 );
not ( n70519 , n69967 );
or ( n70520 , n70222 , n69108 );
nand ( n70521 , n70222 , n2528 );
nand ( n70522 , n70520 , n70521 );
not ( n70523 , n70522 );
nand ( n70524 , n70519 , n70523 );
nand ( n70525 , n70518 , n70524 );
nand ( n70526 , n70517 , n70525 );
nand ( n70527 , n70452 , n70461 );
nand ( n70528 , n70513 , n70515 );
and ( n70529 , n70527 , n70528 );
nand ( n70530 , n70526 , n70529 );
nand ( n70531 , n70464 , n70497 , n70347 , n70530 );
not ( n70532 , n70372 );
and ( n70533 , n70532 , n70283 , n70392 , n70397 );
not ( n70534 , n70489 );
nand ( n70535 , n70425 , n70409 );
not ( n70536 , n70535 );
not ( n70537 , n70438 );
not ( n70538 , n70440 );
nand ( n70539 , n70537 , n70538 );
nand ( n70540 , n70536 , n70539 );
not ( n70541 , n70490 );
nand ( n70542 , n70438 , n70440 );
nand ( n70543 , n70534 , n70540 , n70541 , n70542 );
nand ( n70544 , n70347 , n70497 , n70533 , n70543 );
and ( n70545 , n70384 , n70390 );
not ( n70546 , n70545 );
not ( n70547 , n70397 );
or ( n70548 , n70546 , n70547 );
or ( n70549 , n70394 , n70396 );
nand ( n70550 , n70548 , n70549 );
and ( n70551 , n70550 , n70373 );
nand ( n70552 , n70347 , n70551 );
nand ( n70553 , n70371 , n70531 , n70544 , n70552 );
not ( n70554 , n70553 );
or ( n70555 , n70245 , n70554 );
or ( n70556 , n70553 , n70244 );
nand ( n70557 , n70555 , n70556 );
not ( n70558 , n70188 );
not ( n70559 , n70194 );
nand ( n70560 , n70558 , n70559 );
nand ( n70561 , n70560 , n70195 );
and ( n70562 , n70188 , n70206 );
not ( n70563 , n70188 );
and ( n70564 , n70563 , n70202 );
nor ( n70565 , n70562 , n70564 );
nor ( n70566 , n70561 , n70565 );
not ( n70567 , n70566 );
nor ( n70568 , n70567 , n70183 );
and ( n70569 , n70557 , n70568 );
not ( n70570 , n70565 );
nor ( n70571 , n70570 , n70561 );
not ( n70572 , n70571 );
nor ( n70573 , n70572 , n70183 );
not ( n70574 , n70573 );
not ( n70575 , n70225 );
not ( n70576 , n69641 );
not ( n70577 , n70576 );
or ( n70578 , n70575 , n70577 );
not ( n70579 , n70225 );
nand ( n70580 , n70579 , n69641 );
nand ( n70581 , n70578 , n70580 );
not ( n70582 , n70581 );
and ( n70583 , n69613 , n70238 );
not ( n70584 , n70583 );
nand ( n70585 , n70582 , n70584 );
nand ( n70586 , n70581 , n70583 );
and ( n70587 , n70585 , n70586 );
not ( n70588 , n70587 );
not ( n70589 , n69435 );
not ( n70590 , n70477 );
not ( n70591 , n70590 );
or ( n70592 , n70589 , n70591 );
not ( n70593 , n69435 );
nand ( n70594 , n70593 , n70477 );
nand ( n70595 , n70592 , n70594 );
and ( n70596 , n70432 , n69502 );
nand ( n70597 , n70595 , n70596 );
not ( n70598 , n70597 );
not ( n70599 , n69470 );
not ( n70600 , n70388 );
not ( n70601 , n70600 );
or ( n70602 , n70599 , n70601 );
not ( n70603 , n69470 );
nand ( n70604 , n70603 , n70388 );
nand ( n70605 , n70602 , n70604 );
nand ( n70606 , n70477 , n69435 );
not ( n70607 , n70606 );
nor ( n70608 , n70605 , n70607 );
not ( n70609 , n70608 );
and ( n70610 , n70598 , n70609 );
nand ( n70611 , n70605 , n70607 );
not ( n70612 , n70611 );
nor ( n70613 , n70610 , n70612 );
not ( n70614 , n70595 );
not ( n70615 , n70596 );
nand ( n70616 , n70614 , n70615 );
not ( n70617 , n70608 );
nand ( n70618 , n70616 , n70617 );
nand ( n70619 , n70613 , n70618 );
not ( n70620 , n69543 );
not ( n70621 , n70620 );
not ( n70622 , n70263 );
or ( n70623 , n70621 , n70622 );
not ( n70624 , n70263 );
nand ( n70625 , n70624 , n69543 );
nand ( n70626 , n70623 , n70625 );
not ( n70627 , n70626 );
and ( n70628 , n70378 , n69553 );
not ( n70629 , n70628 );
nand ( n70630 , n70627 , n70629 );
not ( n70631 , n69553 );
not ( n70632 , n70378 );
not ( n70633 , n70632 );
or ( n70634 , n70631 , n70633 );
not ( n70635 , n69553 );
nand ( n70636 , n70378 , n70635 );
nand ( n70637 , n70634 , n70636 );
not ( n70638 , n70637 );
and ( n70639 , n70388 , n69470 );
not ( n70640 , n70639 );
nand ( n70641 , n70638 , n70640 );
nand ( n70642 , n70630 , n70641 );
not ( n70643 , n70273 );
not ( n70644 , n69519 );
not ( n70645 , n70644 );
or ( n70646 , n70643 , n70645 );
not ( n70647 , n70273 );
nand ( n70648 , n69519 , n70647 );
nand ( n70649 , n70646 , n70648 );
not ( n70650 , n70649 );
and ( n70651 , n70253 , n69531 );
not ( n70652 , n70651 );
nand ( n70653 , n70650 , n70652 );
xor ( n70654 , n69531 , n70253 );
not ( n70655 , n70654 );
and ( n70656 , n69543 , n70263 );
not ( n70657 , n70656 );
nand ( n70658 , n70655 , n70657 );
nand ( n70659 , n70653 , n70658 );
nor ( n70660 , n70642 , n70659 );
not ( n70661 , n69576 );
not ( n70662 , n70296 );
not ( n70663 , n70662 );
or ( n70664 , n70661 , n70663 );
not ( n70665 , n69576 );
nand ( n70666 , n70665 , n70296 );
nand ( n70667 , n70664 , n70666 );
nand ( n70668 , n70308 , n69587 );
not ( n70669 , n70668 );
nor ( n70670 , n70667 , n70669 );
not ( n70671 , n70308 );
not ( n70672 , n69587 );
not ( n70673 , n70672 );
or ( n70674 , n70671 , n70673 );
not ( n70675 , n70308 );
nand ( n70676 , n70675 , n69587 );
nand ( n70677 , n70674 , n70676 );
and ( n70678 , n70273 , n69519 );
nor ( n70679 , n70677 , n70678 );
nor ( n70680 , n70670 , n70679 );
not ( n70681 , n70238 );
not ( n70682 , n70681 );
not ( n70683 , n69613 );
or ( n70684 , n70682 , n70683 );
not ( n70685 , n69613 );
nand ( n70686 , n70685 , n70238 );
nand ( n70687 , n70684 , n70686 );
nand ( n70688 , n69599 , n70327 );
not ( n70689 , n70688 );
nor ( n70690 , n70687 , n70689 );
not ( n70691 , n69599 );
not ( n70692 , n70691 );
not ( n70693 , n70327 );
or ( n70694 , n70692 , n70693 );
not ( n70695 , n70327 );
nand ( n70696 , n70695 , n69599 );
nand ( n70697 , n70694 , n70696 );
and ( n70698 , n69576 , n70296 );
nor ( n70699 , n70697 , n70698 );
nor ( n70700 , n70690 , n70699 );
nand ( n70701 , n70619 , n70660 , n70680 , n70700 );
not ( n70702 , n70701 );
not ( n70703 , n70702 );
not ( n70704 , n70459 );
not ( n70705 , n70073 );
not ( n70706 , n70705 );
or ( n70707 , n70704 , n70706 );
not ( n70708 , n70459 );
nand ( n70709 , n70708 , n70073 );
nand ( n70710 , n70707 , n70709 );
not ( n70711 , n70710 );
not ( n70712 , n70053 );
not ( n70713 , n70503 );
nor ( n70714 , n70712 , n70713 );
not ( n70715 , n70714 );
nand ( n70716 , n70711 , n70715 );
not ( n70717 , n70503 );
not ( n70718 , n70053 );
not ( n70719 , n70718 );
or ( n70720 , n70717 , n70719 );
nand ( n70721 , n70053 , n70713 );
nand ( n70722 , n70720 , n70721 );
not ( n70723 , n69967 );
not ( n70724 , n70522 );
nor ( n70725 , n70723 , n70724 );
nand ( n70726 , n70722 , n70725 );
not ( n70727 , n70726 );
nand ( n70728 , n70716 , n70727 );
xor ( n70729 , n69471 , n69451 );
xor ( n70730 , n70729 , n70420 );
and ( n70731 , n70073 , n70459 );
nand ( n70732 , n70730 , n70731 );
nand ( n70733 , n70710 , n70714 );
nand ( n70734 , n70728 , n70732 , n70733 );
not ( n70735 , n69502 );
not ( n70736 , n70432 );
not ( n70737 , n70736 );
or ( n70738 , n70735 , n70737 );
not ( n70739 , n69502 );
nand ( n70740 , n70432 , n70739 );
nand ( n70741 , n70738 , n70740 );
not ( n70742 , n70741 );
and ( n70743 , n70405 , n69487 );
not ( n70744 , n70743 );
nand ( n70745 , n70742 , n70744 );
xor ( n70746 , n69471 , n69451 );
and ( n70747 , n70746 , n70420 );
and ( n70748 , n69471 , n69451 );
or ( n70749 , n70747 , n70748 );
not ( n70750 , n70749 );
not ( n70751 , n69487 );
not ( n70752 , n70405 );
not ( n70753 , n70752 );
or ( n70754 , n70751 , n70753 );
not ( n70755 , n69487 );
nand ( n70756 , n70755 , n70405 );
nand ( n70757 , n70754 , n70756 );
not ( n70758 , n70757 );
nand ( n70759 , n70750 , n70758 );
and ( n70760 , n70745 , n70759 );
or ( n70761 , n70730 , n70731 );
nand ( n70762 , n70734 , n70760 , n70761 );
and ( n70763 , n70749 , n70757 );
not ( n70764 , n70763 );
not ( n70765 , n70745 );
or ( n70766 , n70764 , n70765 );
not ( n70767 , n70744 );
nand ( n70768 , n70767 , n70741 );
nand ( n70769 , n70766 , n70768 );
not ( n70770 , n70613 );
nor ( n70771 , n70769 , n70770 );
nand ( n70772 , n70762 , n70771 );
not ( n70773 , n70772 );
or ( n70774 , n70703 , n70773 );
not ( n70775 , n70697 );
not ( n70776 , n70698 );
nor ( n70777 , n70775 , n70776 );
not ( n70778 , n70777 );
not ( n70779 , n70690 );
not ( n70780 , n70779 );
or ( n70781 , n70778 , n70780 );
nand ( n70782 , n70687 , n70689 );
nand ( n70783 , n70781 , n70782 );
nand ( n70784 , n70677 , n70678 );
or ( n70785 , n70670 , n70784 );
nand ( n70786 , n70667 , n70669 );
nand ( n70787 , n70785 , n70786 );
nor ( n70788 , n70783 , n70787 );
not ( n70789 , n70788 );
nand ( n70790 , n70649 , n70651 );
nand ( n70791 , n70659 , n70790 );
nand ( n70792 , n70654 , n70656 );
nand ( n70793 , n70626 , n70628 );
nand ( n70794 , n70792 , n70790 , n70793 );
not ( n70795 , n70794 );
and ( n70796 , n70637 , n70639 );
nand ( n70797 , n70630 , n70796 );
nand ( n70798 , n70795 , n70797 );
nand ( n70799 , n70791 , n70798 , n70680 );
not ( n70800 , n70799 );
or ( n70801 , n70789 , n70800 );
or ( n70802 , n70783 , n70700 );
nand ( n70803 , n70801 , n70802 );
nand ( n70804 , n70774 , n70803 );
not ( n70805 , n70804 );
not ( n70806 , n70805 );
or ( n70807 , n70588 , n70806 );
nand ( n70808 , n70702 , n70772 );
nand ( n70809 , n70803 , n70808 );
not ( n70810 , n70809 );
or ( n70811 , n70810 , n70587 );
nand ( n70812 , n70807 , n70811 );
not ( n70813 , n70812 );
or ( n70814 , n70574 , n70813 );
not ( n70815 , n70225 );
nor ( n70816 , n70388 , n70432 );
not ( n70817 , n70405 );
not ( n70818 , n70817 );
nor ( n70819 , n70477 , n70818 );
nor ( n70820 , n70327 , n70238 );
nor ( n70821 , n70420 , n70459 );
nand ( n70822 , n70816 , n70819 , n70820 , n70821 );
not ( n70823 , n70822 );
nor ( n70824 , n70263 , n70378 );
not ( n70825 , n70253 );
not ( n70826 , n70273 );
and ( n70827 , n70824 , n70825 , n70826 );
nor ( n70828 , n70296 , n70308 );
not ( n70829 , n70503 );
not ( n70830 , n70829 );
nor ( n70831 , n70830 , n70522 );
nand ( n70832 , n70823 , n70827 , n70828 , n70831 );
not ( n70833 , n70832 );
not ( n70834 , n70833 );
or ( n70835 , n70815 , n70834 );
or ( n70836 , n70833 , n70225 );
nand ( n70837 , n70835 , n70836 );
nor ( n70838 , n70188 , n70194 );
nand ( n70839 , n70838 , n70207 );
nor ( n70840 , n70183 , n70839 );
nand ( n70841 , n70837 , n70840 );
not ( n70842 , n70183 );
not ( n70843 , n70194 );
not ( n70844 , n70202 );
nor ( n70845 , n70844 , n70188 );
nand ( n70846 , n70843 , n70845 );
not ( n70847 , n70846 );
nand ( n70848 , n70842 , n70847 );
not ( n70849 , n70848 );
nand ( n70850 , n70849 , n70225 );
not ( n70851 , n70845 );
nor ( n70852 , n70202 , n70206 );
not ( n70853 , n70852 );
nand ( n70854 , n70561 , n70851 , n70853 );
not ( n70855 , n70854 );
not ( n70856 , n70164 );
or ( n70857 , n70855 , n70856 );
or ( n70858 , n70195 , n70207 );
not ( n70859 , n70139 );
not ( n70860 , n70859 );
nand ( n70861 , n70136 , n70860 );
not ( n70862 , n70861 );
not ( n70863 , n70147 );
nand ( n70864 , n70858 , n70862 , n70863 );
not ( n70865 , n70206 );
nor ( n70866 , n70202 , n70865 );
and ( n70867 , n70838 , n70866 );
nor ( n70868 , n70867 , n70180 );
nor ( n70869 , n70864 , n70868 );
nand ( n70870 , n70857 , n70869 );
and ( n70871 , n70870 , n2697 );
not ( n70872 , n70560 );
nand ( n70873 , n70866 , n70139 );
not ( n70874 , n70873 );
nand ( n70875 , n70136 , n70872 , n70874 , n70863 );
not ( n70876 , n70875 );
not ( n70877 , n3356 );
nand ( n70878 , n3304 , n3344 );
nor ( n70879 , n70877 , n70878 );
nand ( n70880 , n70879 , n3288 );
not ( n70881 , n3324 );
nor ( n70882 , n70880 , n70881 );
nand ( n70883 , n70882 , n69549 );
not ( n70884 , n69537 );
nor ( n70885 , n70883 , n70884 );
nand ( n70886 , n70885 , n69520 );
not ( n70887 , n69512 );
nor ( n70888 , n70886 , n70887 );
and ( n70889 , n70888 , n3442 );
nand ( n70890 , n70889 , n69567 );
not ( n70891 , n3454 );
nor ( n70892 , n70890 , n70891 );
nand ( n70893 , n70892 , n69603 );
not ( n70894 , n69639 );
and ( n70895 , n70893 , n70894 );
not ( n70896 , n70893 );
and ( n70897 , n70896 , n69639 );
nor ( n70898 , n70895 , n70897 );
and ( n70899 , n70876 , n70898 );
nor ( n70900 , n70871 , n70899 );
and ( n70901 , n70841 , n70850 , n70900 );
nand ( n70902 , n70814 , n70901 );
nor ( n70903 , n70569 , n70902 );
nand ( n70904 , n70211 , n70903 );
buf ( n70905 , n70904 );
buf ( n70906 , 1'b0 );
not ( n70907 , n68838 );
buf ( n4769 , n70907 );
buf ( n4770 , n68634 );
not ( n70910 , n69358 );
not ( n70911 , n70013 );
nand ( n70912 , n69969 , n70092 );
not ( n70913 , n70912 );
nand ( n70914 , n70913 , n70007 );
not ( n70915 , n70914 );
or ( n70916 , n70911 , n70915 );
or ( n70917 , n70914 , n70013 );
nand ( n70918 , n70916 , n70917 );
not ( n70919 , n70918 );
or ( n70920 , n70910 , n70919 );
nand ( n70921 , n70082 , n69359 );
nand ( n70922 , n70920 , n70921 );
not ( n70923 , n70195 );
and ( n70924 , n70922 , n70923 );
not ( n70925 , n70206 );
not ( n70926 , n70188 );
or ( n70927 , n70925 , n70926 );
or ( n70928 , n70872 , n70851 );
nand ( n70929 , n70927 , n70928 );
not ( n70930 , n70929 );
not ( n70931 , n70930 );
not ( n70932 , n70931 );
nand ( n70933 , n70397 , n70549 );
not ( n70934 , n70933 );
not ( n70935 , n70392 );
not ( n70936 , n70442 );
nor ( n70937 , n70496 , n70936 );
not ( n70938 , n70937 );
not ( n70939 , n70463 );
not ( n70940 , n70526 );
not ( n70941 , n70940 );
or ( n70942 , n70939 , n70941 );
not ( n70943 , n70528 );
and ( n70944 , n70463 , n70943 );
not ( n70945 , n70527 );
nor ( n70946 , n70944 , n70945 );
nand ( n70947 , n70942 , n70946 );
not ( n70948 , n70947 );
or ( n70949 , n70938 , n70948 );
nand ( n70950 , n70540 , n70542 );
not ( n70951 , n70950 );
not ( n70952 , n70496 );
not ( n70953 , n70952 );
or ( n70954 , n70951 , n70953 );
nand ( n70955 , n70954 , n70491 );
not ( n70956 , n70955 );
nand ( n70957 , n70949 , n70956 );
not ( n70958 , n70957 );
or ( n70959 , n70935 , n70958 );
not ( n70960 , n70545 );
nand ( n70961 , n70959 , n70960 );
not ( n70962 , n70961 );
or ( n70963 , n70934 , n70962 );
or ( n70964 , n70961 , n70933 );
nand ( n70965 , n70963 , n70964 );
not ( n70966 , n70965 );
or ( n70967 , n70932 , n70966 );
nand ( n70968 , n70630 , n70793 );
not ( n70969 , n70968 );
not ( n70970 , n70641 );
not ( n70971 , n70760 );
nor ( n70972 , n70971 , n70618 );
not ( n70973 , n70972 );
not ( n70974 , n70728 );
nand ( n70975 , n70974 , n70761 );
not ( n70976 , n70733 );
nand ( n70977 , n70761 , n70976 );
nand ( n70978 , n70975 , n70977 , n70732 );
not ( n70979 , n70978 );
or ( n70980 , n70973 , n70979 );
not ( n70981 , n70618 );
and ( n70982 , n70769 , n70981 );
nor ( n70983 , n70982 , n70770 );
nand ( n70984 , n70980 , n70983 );
not ( n70985 , n70984 );
or ( n70986 , n70970 , n70985 );
not ( n70987 , n70796 );
nand ( n70988 , n70986 , n70987 );
not ( n70989 , n70988 );
or ( n70990 , n70969 , n70989 );
or ( n70991 , n70988 , n70968 );
nand ( n70992 , n70990 , n70991 );
and ( n70993 , n70992 , n70571 );
not ( n70994 , n70852 );
nor ( n70995 , n70994 , n70560 );
not ( n70996 , n70995 );
not ( n70997 , n70263 );
not ( n70998 , n70997 );
not ( n70999 , n70378 );
and ( n71000 , n70831 , n70821 );
and ( n71001 , n70819 , n70816 );
nand ( n71002 , n71000 , n71001 );
not ( n71003 , n71002 );
nand ( n71004 , n70999 , n71003 );
not ( n71005 , n71004 );
or ( n71006 , n70998 , n71005 );
or ( n71007 , n71004 , n70997 );
nand ( n71008 , n71006 , n71007 );
not ( n71009 , n71008 );
or ( n71010 , n70996 , n71009 );
nand ( n71011 , n70847 , n70263 );
nand ( n71012 , n71010 , n71011 );
nor ( n71013 , n70993 , n71012 );
nand ( n71014 , n70967 , n71013 );
nor ( n71015 , n70924 , n71014 );
nand ( n71016 , n70148 , n70164 , n70181 , n70854 );
or ( n71017 , n71015 , n71016 );
nand ( n71018 , n71016 , n69535 );
nand ( n71019 , n71017 , n71018 );
buf ( n4881 , n71019 );
buf ( n71021 , 1'b0 );
not ( n71022 , n68838 );
buf ( n4884 , n71022 );
buf ( n4885 , n68634 );
not ( n71025 , n71016 );
not ( n71026 , n69800 );
or ( n71027 , n71025 , n71026 );
not ( n71028 , n69358 );
nor ( n71029 , n69823 , n69826 );
not ( n71030 , n71029 );
not ( n71031 , n71030 );
nand ( n71032 , n71031 , n69627 );
not ( n71033 , n69871 );
and ( n71034 , n71032 , n71033 );
not ( n71035 , n71032 );
and ( n71036 , n71035 , n69871 );
nor ( n71037 , n71034 , n71036 );
not ( n71038 , n71037 );
nand ( n71039 , n69983 , n69660 );
nor ( n71040 , n70099 , n71039 );
nand ( n71041 , n69971 , n71040 );
nand ( n71042 , n69627 , n69827 );
not ( n71043 , n69822 );
and ( n71044 , n71042 , n71043 );
not ( n71045 , n71042 );
and ( n71046 , n71045 , n69822 );
nor ( n71047 , n71044 , n71046 );
not ( n71048 , n71047 );
nor ( n71049 , n71041 , n71048 );
not ( n71050 , n69804 );
not ( n71051 , n69827 );
nor ( n71052 , n71051 , n71043 );
nand ( n71053 , n69627 , n71052 );
not ( n71054 , n71053 );
or ( n71055 , n71050 , n71054 );
nand ( n71056 , n69627 , n71052 );
or ( n71057 , n71056 , n69804 );
nand ( n71058 , n71055 , n71057 );
nand ( n71059 , n71049 , n71058 );
not ( n71060 , n71059 );
or ( n71061 , n71038 , n71060 );
or ( n71062 , n71059 , n71037 );
nand ( n71063 , n71061 , n71062 );
not ( n71064 , n71063 );
or ( n71065 , n71028 , n71064 );
nand ( n71066 , n71047 , n69359 );
nand ( n71067 , n71065 , n71066 );
and ( n71068 , n71067 , n70923 );
not ( n71069 , n69176 );
not ( n71070 , n70222 );
not ( n71071 , n71070 );
or ( n71072 , n71069 , n71071 );
nand ( n71073 , n70222 , n68650 );
nand ( n71074 , n71072 , n71073 );
not ( n71075 , n71074 );
not ( n71076 , n71075 );
not ( n71077 , n69655 );
not ( n71078 , n71077 );
or ( n71079 , n71076 , n71078 );
nand ( n71080 , n69655 , n71074 );
nand ( n71081 , n71079 , n71080 );
nand ( n71082 , n70229 , n69641 );
not ( n71083 , n71082 );
nor ( n71084 , n71081 , n71083 );
nor ( n71085 , n71084 , n70241 );
not ( n71086 , n71085 );
not ( n71087 , n69822 );
not ( n71088 , n69157 );
not ( n71089 , n71070 );
or ( n71090 , n71088 , n71089 );
nand ( n71091 , n70222 , n68649 );
nand ( n71092 , n71090 , n71091 );
not ( n71093 , n71092 );
or ( n71094 , n71087 , n71093 );
not ( n71095 , n71092 );
not ( n71096 , n69822 );
nand ( n71097 , n71095 , n71096 );
nand ( n71098 , n71094 , n71097 );
and ( n71099 , n71075 , n69655 );
nor ( n71100 , n71098 , n71099 );
nor ( n71101 , n71086 , n71100 );
not ( n71102 , n71101 );
not ( n71103 , n70553 );
or ( n71104 , n71102 , n71103 );
not ( n71105 , n71100 );
not ( n71106 , n71105 );
or ( n71107 , n70243 , n71084 );
nand ( n71108 , n71081 , n71083 );
nand ( n71109 , n71107 , n71108 );
not ( n71110 , n71109 );
or ( n71111 , n71106 , n71110 );
nand ( n71112 , n71098 , n71099 );
nand ( n71113 , n71111 , n71112 );
not ( n71114 , n71113 );
nand ( n71115 , n71104 , n71114 );
not ( n71116 , n69804 );
not ( n71117 , n70222 );
not ( n71118 , n69241 );
and ( n71119 , n71117 , n71118 );
and ( n71120 , n70222 , n2509 );
nor ( n71121 , n71119 , n71120 );
not ( n71122 , n71121 );
not ( n71123 , n71122 );
or ( n71124 , n71116 , n71123 );
not ( n71125 , n71122 );
not ( n71126 , n69804 );
nand ( n71127 , n71125 , n71126 );
nand ( n71128 , n71124 , n71127 );
not ( n71129 , n69822 );
nor ( n71130 , n71129 , n71092 );
nor ( n71131 , n71128 , n71130 );
and ( n71132 , n71128 , n71130 );
or ( n71133 , n71131 , n71132 );
xnor ( n71134 , n71115 , n71133 );
nand ( n71135 , n71134 , n70929 );
not ( n71136 , n71122 );
not ( n71137 , n71136 );
not ( n71138 , n69804 );
or ( n71139 , n71137 , n71138 );
not ( n71140 , n69804 );
nand ( n71141 , n71140 , n71122 );
nand ( n71142 , n71139 , n71141 );
nand ( n71143 , n71092 , n69822 );
not ( n71144 , n71143 );
and ( n71145 , n71142 , n71144 );
nor ( n71146 , n71142 , n71144 );
or ( n71147 , n71145 , n71146 );
not ( n71148 , n71147 );
not ( n71149 , n69655 );
not ( n71150 , n71074 );
not ( n71151 , n71150 );
or ( n71152 , n71149 , n71151 );
not ( n71153 , n69655 );
nand ( n71154 , n71153 , n71074 );
nand ( n71155 , n71152 , n71154 );
nand ( n71156 , n69641 , n70225 );
not ( n71157 , n71156 );
nor ( n71158 , n71155 , n71157 );
not ( n71159 , n71158 );
nand ( n71160 , n71159 , n70585 );
not ( n71161 , n69822 );
not ( n71162 , n71092 );
not ( n71163 , n71162 );
or ( n71164 , n71161 , n71163 );
not ( n71165 , n69822 );
nand ( n71166 , n71092 , n71165 );
nand ( n71167 , n71164 , n71166 );
and ( n71168 , n69655 , n71074 );
nor ( n71169 , n71167 , n71168 );
nor ( n71170 , n71160 , n71169 );
not ( n71171 , n71170 );
not ( n71172 , n70804 );
or ( n71173 , n71171 , n71172 );
not ( n71174 , n71169 );
not ( n71175 , n71174 );
or ( n71176 , n71158 , n70586 );
nand ( n71177 , n71155 , n71157 );
nand ( n71178 , n71176 , n71177 );
not ( n71179 , n71178 );
or ( n71180 , n71175 , n71179 );
nand ( n71181 , n71167 , n71168 );
nand ( n71182 , n71180 , n71181 );
not ( n71183 , n71182 );
nand ( n71184 , n71173 , n71183 );
not ( n71185 , n71184 );
or ( n71186 , n71148 , n71185 );
or ( n71187 , n71184 , n71147 );
nand ( n71188 , n71186 , n71187 );
and ( n71189 , n71188 , n70571 );
not ( n71190 , n70995 );
not ( n71191 , n71122 );
not ( n71192 , n70225 );
not ( n71193 , n71074 );
nand ( n71194 , n71192 , n71193 );
or ( n71195 , n71194 , n71092 );
nor ( n71196 , n70832 , n71195 );
not ( n71197 , n71196 );
or ( n71198 , n71191 , n71197 );
or ( n71199 , n71196 , n71122 );
nand ( n71200 , n71198 , n71199 );
not ( n71201 , n71200 );
or ( n71202 , n71190 , n71201 );
nand ( n71203 , n70847 , n71122 );
nand ( n71204 , n71202 , n71203 );
nor ( n71205 , n71189 , n71204 );
nand ( n71206 , n71135 , n71205 );
nor ( n71207 , n71068 , n71206 );
or ( n71208 , n71207 , n71016 );
nand ( n71209 , n71027 , n71208 );
buf ( n5071 , n71209 );
buf ( n5072 , 1'b0 );
not ( n71212 , n68838 );
buf ( n5074 , n71212 );
buf ( n5075 , n68634 );
not ( n71215 , n69358 );
not ( n71216 , n71058 );
not ( n71217 , n71216 );
not ( n71218 , n71049 );
or ( n71219 , n71217 , n71218 );
or ( n71220 , n71049 , n71216 );
nand ( n71221 , n71219 , n71220 );
not ( n71222 , n71221 );
or ( n71223 , n71215 , n71222 );
nand ( n71224 , n69660 , n69359 );
nand ( n71225 , n71223 , n71224 );
and ( n71226 , n71225 , n70923 );
not ( n71227 , n71085 );
not ( n71228 , n70553 );
or ( n71229 , n71227 , n71228 );
not ( n71230 , n71109 );
nand ( n71231 , n71229 , n71230 );
nand ( n71232 , n71105 , n71112 );
xnor ( n71233 , n71231 , n71232 );
not ( n71234 , n71233 );
not ( n71235 , n70929 );
or ( n71236 , n71234 , n71235 );
nand ( n71237 , n71174 , n71181 );
not ( n71238 , n71237 );
not ( n71239 , n71160 );
not ( n71240 , n71239 );
not ( n71241 , n70804 );
or ( n71242 , n71240 , n71241 );
not ( n71243 , n71178 );
nand ( n71244 , n71242 , n71243 );
not ( n71245 , n71244 );
or ( n71246 , n71238 , n71245 );
or ( n71247 , n71244 , n71237 );
nand ( n71248 , n71246 , n71247 );
and ( n71249 , n71248 , n70571 );
not ( n71250 , n70995 );
not ( n71251 , n71092 );
nor ( n71252 , n70832 , n71194 );
not ( n71253 , n71252 );
or ( n71254 , n71251 , n71253 );
or ( n71255 , n71252 , n71092 );
nand ( n71256 , n71254 , n71255 );
not ( n71257 , n71256 );
or ( n71258 , n71250 , n71257 );
nand ( n71259 , n70847 , n71092 );
nand ( n71260 , n71258 , n71259 );
nor ( n71261 , n71249 , n71260 );
nand ( n71262 , n71236 , n71261 );
nor ( n71263 , n71226 , n71262 );
or ( n71264 , n71263 , n71016 );
nand ( n71265 , n71016 , n69810 );
nand ( n71266 , n71264 , n71265 );
buf ( n5128 , n71266 );
buf ( n71268 , 1'b0 );
not ( n71269 , n68838 );
buf ( n71270 , n71269 );
buf ( n5132 , n68634 );
not ( n71272 , n69358 );
and ( n71273 , n71272 , n69977 );
not ( n71274 , n71272 );
not ( n71275 , n71047 );
not ( n71276 , n71041 );
or ( n71277 , n71275 , n71276 );
or ( n71278 , n71041 , n71047 );
nand ( n71279 , n71277 , n71278 );
and ( n71280 , n71274 , n71279 );
nor ( n71281 , n71273 , n71280 );
not ( n71282 , n71281 );
and ( n71283 , n71282 , n70923 );
not ( n71284 , n70929 );
not ( n71285 , n70242 );
not ( n71286 , n70553 );
or ( n71287 , n71285 , n71286 );
nand ( n71288 , n71287 , n70243 );
not ( n71289 , n71084 );
nand ( n71290 , n71289 , n71108 );
xnor ( n71291 , n71288 , n71290 );
not ( n71292 , n71291 );
or ( n71293 , n71284 , n71292 );
not ( n71294 , n71158 );
nand ( n71295 , n71294 , n71177 );
not ( n71296 , n71295 );
not ( n71297 , n70585 );
not ( n71298 , n70804 );
or ( n71299 , n71297 , n71298 );
nand ( n71300 , n71299 , n70586 );
not ( n71301 , n71300 );
or ( n71302 , n71296 , n71301 );
or ( n71303 , n71300 , n71295 );
nand ( n71304 , n71302 , n71303 );
and ( n71305 , n71304 , n70571 );
not ( n71306 , n70995 );
not ( n71307 , n71074 );
nor ( n71308 , n70832 , n70225 );
not ( n71309 , n71308 );
or ( n71310 , n71307 , n71309 );
or ( n71311 , n71308 , n71074 );
nand ( n71312 , n71310 , n71311 );
not ( n71313 , n71312 );
or ( n71314 , n71306 , n71313 );
nand ( n71315 , n70847 , n71074 );
nand ( n71316 , n71314 , n71315 );
nor ( n71317 , n71305 , n71316 );
nand ( n71318 , n71293 , n71317 );
nor ( n71319 , n71283 , n71318 );
or ( n71320 , n71319 , n71016 );
nand ( n71321 , n71016 , n3510 );
nand ( n71322 , n71320 , n71321 );
buf ( n71323 , n71322 );
buf ( n71324 , 1'b0 );
not ( n71325 , n68838 );
buf ( n71326 , n71325 );
buf ( n71327 , n68634 );
not ( n71328 , n70109 );
and ( n71329 , n71328 , n70196 );
not ( n71330 , n70931 );
not ( n71331 , n70557 );
or ( n71332 , n71330 , n71331 );
and ( n71333 , n70812 , n70571 );
not ( n71334 , n70995 );
not ( n71335 , n70837 );
or ( n71336 , n71334 , n71335 );
nand ( n71337 , n70225 , n70847 );
nand ( n71338 , n71336 , n71337 );
nor ( n71339 , n71333 , n71338 );
nand ( n71340 , n71332 , n71339 );
nor ( n71341 , n71329 , n71340 );
or ( n71342 , n71341 , n71016 );
not ( n71343 , n71016 );
not ( n71344 , n71343 );
nand ( n71345 , n71344 , n3498 );
nand ( n71346 , n71342 , n71345 );
buf ( n71347 , n71346 );
buf ( n71348 , 1'b0 );
not ( n71349 , n68838 );
buf ( n71350 , n71349 );
buf ( n71351 , n68634 );
not ( n71352 , n69358 );
not ( n71353 , n69978 );
not ( n71354 , n71353 );
nor ( n71355 , n70101 , n69982 );
nand ( n71356 , n69969 , n71355 );
not ( n71357 , n71356 );
or ( n71358 , n71354 , n71357 );
or ( n71359 , n71356 , n71353 );
nand ( n71360 , n71358 , n71359 );
not ( n71361 , n71360 );
or ( n71362 , n71352 , n71361 );
nand ( n71363 , n69981 , n71272 );
nand ( n71364 , n71362 , n71363 );
and ( n71365 , n71364 , n70196 );
not ( n71366 , n70931 );
not ( n71367 , n70345 );
nand ( n71368 , n71367 , n70365 );
not ( n71369 , n71368 );
not ( n71370 , n70336 );
nand ( n71371 , n70321 , n71370 );
not ( n71372 , n70533 );
nor ( n71373 , n71371 , n71372 );
not ( n71374 , n71373 );
not ( n71375 , n70957 );
or ( n71376 , n71374 , n71375 );
nor ( n71377 , n70287 , n70551 );
not ( n71378 , n71377 );
not ( n71379 , n71371 );
and ( n71380 , n71378 , n71379 );
not ( n71381 , n71370 );
not ( n71382 , n70358 );
or ( n71383 , n71381 , n71382 );
nand ( n71384 , n71383 , n70362 );
nor ( n71385 , n71380 , n71384 );
nand ( n71386 , n71376 , n71385 );
not ( n71387 , n71386 );
or ( n71388 , n71369 , n71387 );
or ( n71389 , n71386 , n71368 );
nand ( n71390 , n71388 , n71389 );
not ( n71391 , n71390 );
or ( n71392 , n71366 , n71391 );
nand ( n71393 , n70779 , n70782 );
not ( n71394 , n71393 );
not ( n71395 , n70699 );
nand ( n71396 , n70680 , n71395 );
not ( n71397 , n70660 );
nor ( n71398 , n71396 , n71397 );
not ( n71399 , n71398 );
not ( n71400 , n70984 );
or ( n71401 , n71399 , n71400 );
nand ( n71402 , n70798 , n70791 );
not ( n71403 , n71402 );
not ( n71404 , n71396 );
and ( n71405 , n71403 , n71404 );
not ( n71406 , n71395 );
not ( n71407 , n70787 );
or ( n71408 , n71406 , n71407 );
not ( n71409 , n70777 );
nand ( n71410 , n71408 , n71409 );
nor ( n71411 , n71405 , n71410 );
nand ( n71412 , n71401 , n71411 );
not ( n71413 , n71412 );
or ( n71414 , n71394 , n71413 );
or ( n71415 , n71412 , n71393 );
nand ( n71416 , n71414 , n71415 );
and ( n71417 , n71416 , n70571 );
not ( n71418 , n70995 );
not ( n71419 , n70238 );
not ( n71420 , n71419 );
not ( n71421 , n70327 );
nand ( n71422 , n70827 , n70828 , n71421 );
not ( n71423 , n71422 );
nand ( n71424 , n71423 , n71003 );
not ( n71425 , n71424 );
or ( n71426 , n71420 , n71425 );
or ( n71427 , n71424 , n71419 );
nand ( n71428 , n71426 , n71427 );
not ( n71429 , n71428 );
or ( n71430 , n71418 , n71429 );
nand ( n71431 , n70238 , n70847 );
nand ( n71432 , n71430 , n71431 );
nor ( n71433 , n71417 , n71432 );
nand ( n71434 , n71392 , n71433 );
nor ( n71435 , n71365 , n71434 );
or ( n71436 , n71435 , n71016 );
nand ( n71437 , n71016 , n69607 );
nand ( n71438 , n71436 , n71437 );
buf ( n5300 , n71438 );
buf ( n71440 , 1'b0 );
not ( n71441 , n68838 );
buf ( n71442 , n71441 );
buf ( n5304 , n68634 );
not ( n71444 , n69358 );
not ( n71445 , n69618 );
not ( n71446 , n71445 );
nand ( n71447 , n69969 , n70100 );
not ( n71448 , n69981 );
nor ( n71449 , n71447 , n71448 );
not ( n71450 , n71449 );
or ( n71451 , n71446 , n71450 );
or ( n71452 , n71449 , n71445 );
nand ( n71453 , n71451 , n71452 );
not ( n71454 , n71453 );
or ( n71455 , n71444 , n71454 );
nand ( n71456 , n70098 , n69359 );
nand ( n71457 , n71455 , n71456 );
and ( n71458 , n71457 , n70923 );
not ( n71459 , n70929 );
nand ( n71460 , n71370 , n70362 );
not ( n71461 , n71460 );
not ( n71462 , n70321 );
nor ( n71463 , n71372 , n71462 );
not ( n71464 , n71463 );
not ( n71465 , n70957 );
or ( n71466 , n71464 , n71465 );
or ( n71467 , n71377 , n71462 );
not ( n71468 , n70358 );
nand ( n71469 , n71467 , n71468 );
not ( n71470 , n71469 );
nand ( n71471 , n71466 , n71470 );
not ( n71472 , n71471 );
or ( n71473 , n71461 , n71472 );
or ( n71474 , n71471 , n71460 );
nand ( n71475 , n71473 , n71474 );
not ( n71476 , n71475 );
or ( n71477 , n71459 , n71476 );
nand ( n71478 , n71395 , n71409 );
not ( n71479 , n71478 );
not ( n71480 , n70680 );
nor ( n71481 , n71480 , n71397 );
not ( n71482 , n71481 );
not ( n71483 , n70984 );
or ( n71484 , n71482 , n71483 );
not ( n71485 , n70799 );
nor ( n71486 , n71485 , n70787 );
nand ( n71487 , n71484 , n71486 );
not ( n71488 , n71487 );
or ( n71489 , n71479 , n71488 );
or ( n71490 , n71487 , n71478 );
nand ( n71491 , n71489 , n71490 );
and ( n71492 , n71491 , n70571 );
not ( n71493 , n70995 );
not ( n71494 , n71421 );
nand ( n71495 , n70827 , n70828 );
not ( n71496 , n71495 );
nand ( n71497 , n71496 , n71003 );
not ( n71498 , n71497 );
or ( n71499 , n71494 , n71498 );
or ( n71500 , n71497 , n71421 );
nand ( n71501 , n71499 , n71500 );
not ( n71502 , n71501 );
or ( n71503 , n71493 , n71502 );
nand ( n71504 , n70327 , n70847 );
nand ( n71505 , n71503 , n71504 );
nor ( n71506 , n71492 , n71505 );
nand ( n71507 , n71477 , n71506 );
nor ( n71508 , n71458 , n71507 );
or ( n71509 , n71508 , n71016 );
nand ( n71510 , n71016 , n69591 );
nand ( n71511 , n71509 , n71510 );
buf ( n71512 , n71511 );
buf ( n5374 , 1'b0 );
not ( n71514 , n68838 );
buf ( n71515 , n71514 );
buf ( n71516 , n68634 );
not ( n71517 , n69358 );
not ( n71518 , n70098 );
not ( n71519 , n70015 );
not ( n71520 , n70001 );
and ( n71521 , n70092 , n71519 , n71520 );
nand ( n71522 , n69971 , n71521 );
not ( n71523 , n71522 );
or ( n71524 , n71518 , n71523 );
or ( n71525 , n71522 , n70098 );
nand ( n71526 , n71524 , n71525 );
not ( n71527 , n71526 );
or ( n71528 , n71517 , n71527 );
not ( n71529 , n70000 );
not ( n71530 , n71529 );
nand ( n71531 , n71530 , n69359 );
nand ( n71532 , n71528 , n71531 );
and ( n71533 , n71532 , n70923 );
not ( n71534 , n70931 );
not ( n71535 , n70320 );
nand ( n71536 , n71535 , n70351 );
not ( n71537 , n71536 );
not ( n71538 , n70533 );
not ( n71539 , n70957 );
or ( n71540 , n71538 , n71539 );
nand ( n71541 , n71540 , n71377 );
not ( n71542 , n71541 );
or ( n71543 , n71537 , n71542 );
or ( n71544 , n71541 , n71536 );
nand ( n71545 , n71543 , n71544 );
not ( n71546 , n71545 );
or ( n71547 , n71534 , n71546 );
not ( n71548 , n70679 );
nand ( n71549 , n71548 , n70784 );
not ( n71550 , n71549 );
not ( n71551 , n70660 );
not ( n71552 , n70984 );
or ( n71553 , n71551 , n71552 );
nand ( n71554 , n71553 , n71402 );
not ( n71555 , n71554 );
or ( n71556 , n71550 , n71555 );
or ( n71557 , n71554 , n71549 );
nand ( n71558 , n71556 , n71557 );
and ( n71559 , n71558 , n70571 );
not ( n71560 , n70995 );
not ( n71561 , n70308 );
not ( n71562 , n71561 );
nand ( n71563 , n71003 , n70827 );
not ( n71564 , n71563 );
or ( n71565 , n71562 , n71564 );
or ( n71566 , n71563 , n71561 );
nand ( n71567 , n71565 , n71566 );
not ( n71568 , n71567 );
or ( n71569 , n71560 , n71568 );
nand ( n71570 , n70308 , n70847 );
nand ( n71571 , n71569 , n71570 );
nor ( n71572 , n71559 , n71571 );
nand ( n71573 , n71547 , n71572 );
nor ( n71574 , n71533 , n71573 );
or ( n71575 , n71574 , n71016 );
nand ( n71576 , n71016 , n69579 );
nand ( n71577 , n71575 , n71576 );
buf ( n5439 , n71577 );
buf ( n5440 , 1'b0 );
not ( n71580 , n68838 );
buf ( n71581 , n71580 );
buf ( n71582 , n68634 );
not ( n71583 , n69358 );
not ( n71584 , n69990 );
not ( n71585 , n71584 );
not ( n71586 , n70091 );
and ( n71587 , n71586 , n70014 );
nand ( n71588 , n69969 , n71587 );
not ( n71589 , n70000 );
nor ( n71590 , n71588 , n71589 );
not ( n71591 , n71590 );
or ( n71592 , n71585 , n71591 );
or ( n71593 , n71590 , n71584 );
nand ( n71594 , n71592 , n71593 );
not ( n71595 , n71594 );
or ( n71596 , n71583 , n71595 );
nand ( n71597 , n70013 , n69359 );
nand ( n71598 , n71596 , n71597 );
and ( n71599 , n71598 , n70196 );
not ( n71600 , n70931 );
nand ( n71601 , n70283 , n70286 );
not ( n71602 , n71601 );
not ( n71603 , n70398 );
nor ( n71604 , n71603 , n70372 );
not ( n71605 , n71604 );
not ( n71606 , n70957 );
or ( n71607 , n71605 , n71606 );
not ( n71608 , n70532 );
not ( n71609 , n70550 );
or ( n71610 , n71608 , n71609 );
not ( n71611 , n70266 );
nand ( n71612 , n71610 , n71611 );
not ( n71613 , n71612 );
nand ( n71614 , n71607 , n71613 );
not ( n71615 , n71614 );
or ( n71616 , n71602 , n71615 );
or ( n71617 , n71614 , n71601 );
nand ( n71618 , n71616 , n71617 );
not ( n71619 , n71618 );
or ( n71620 , n71600 , n71619 );
nand ( n71621 , n70653 , n70790 );
not ( n71622 , n71621 );
not ( n71623 , n70658 );
nor ( n71624 , n71623 , n70642 );
not ( n71625 , n71624 );
not ( n71626 , n70984 );
or ( n71627 , n71625 , n71626 );
not ( n71628 , n70658 );
nand ( n71629 , n70797 , n70793 );
not ( n71630 , n71629 );
or ( n71631 , n71628 , n71630 );
nand ( n71632 , n71631 , n70792 );
not ( n71633 , n71632 );
nand ( n71634 , n71627 , n71633 );
not ( n71635 , n71634 );
or ( n71636 , n71622 , n71635 );
or ( n71637 , n71634 , n71621 );
nand ( n71638 , n71636 , n71637 );
and ( n71639 , n71638 , n70571 );
not ( n71640 , n70995 );
not ( n71641 , n70826 );
and ( n71642 , n70824 , n70825 );
nand ( n71643 , n71003 , n71642 );
not ( n71644 , n71643 );
or ( n71645 , n71641 , n71644 );
or ( n71646 , n71643 , n70826 );
nand ( n71647 , n71645 , n71646 );
not ( n71648 , n71647 );
or ( n71649 , n71640 , n71648 );
nand ( n71650 , n70273 , n70847 );
nand ( n71651 , n71649 , n71650 );
nor ( n71652 , n71639 , n71651 );
nand ( n71653 , n71620 , n71652 );
nor ( n71654 , n71599 , n71653 );
or ( n71655 , n71654 , n71016 );
nand ( n71656 , n71016 , n69509 );
nand ( n71657 , n71655 , n71656 );
buf ( n71658 , n71657 );
buf ( n71659 , 1'b0 );
not ( n71660 , n68838 );
buf ( n71661 , n71660 );
buf ( n71662 , n68634 );
not ( n71663 , n69358 );
not ( n71664 , n70000 );
not ( n71665 , n71588 );
or ( n71666 , n71664 , n71665 );
or ( n71667 , n71588 , n70000 );
nand ( n71668 , n71666 , n71667 );
not ( n71669 , n71668 );
or ( n71670 , n71663 , n71669 );
nand ( n71671 , n70007 , n69359 );
nand ( n71672 , n71670 , n71671 );
and ( n71673 , n71672 , n70196 );
not ( n71674 , n70929 );
nand ( n71675 , n70532 , n71611 );
not ( n71676 , n71675 );
not ( n71677 , n70398 );
not ( n71678 , n70957 );
or ( n71679 , n71677 , n71678 );
not ( n71680 , n70550 );
nand ( n71681 , n71679 , n71680 );
not ( n71682 , n71681 );
or ( n71683 , n71676 , n71682 );
or ( n71684 , n71681 , n71675 );
nand ( n71685 , n71683 , n71684 );
not ( n71686 , n71685 );
or ( n71687 , n71674 , n71686 );
nand ( n71688 , n70658 , n70792 );
not ( n71689 , n71688 );
not ( n71690 , n70642 );
not ( n71691 , n71690 );
not ( n71692 , n70984 );
or ( n71693 , n71691 , n71692 );
not ( n71694 , n71629 );
nand ( n71695 , n71693 , n71694 );
not ( n71696 , n71695 );
or ( n71697 , n71689 , n71696 );
or ( n71698 , n71695 , n71688 );
nand ( n71699 , n71697 , n71698 );
and ( n71700 , n71699 , n70571 );
not ( n71701 , n70995 );
not ( n71702 , n70825 );
nand ( n71703 , n71003 , n70824 );
not ( n71704 , n71703 );
or ( n71705 , n71702 , n71704 );
or ( n71706 , n71703 , n70825 );
nand ( n71707 , n71705 , n71706 );
not ( n71708 , n71707 );
or ( n71709 , n71701 , n71708 );
nand ( n71710 , n70253 , n70847 );
nand ( n71711 , n71709 , n71710 );
nor ( n71712 , n71700 , n71711 );
nand ( n71713 , n71687 , n71712 );
nor ( n71714 , n71673 , n71713 );
or ( n71715 , n71714 , n71016 );
nand ( n71716 , n71016 , n69524 );
nand ( n71717 , n71715 , n71716 );
buf ( n71718 , n71717 );
buf ( n71719 , 1'b0 );
not ( n71720 , n68838 );
buf ( n5582 , n71720 );
buf ( n71722 , n68634 );
nand ( n71723 , n70146 , n70860 );
nor ( n71724 , n70136 , n71723 );
not ( n71725 , n71724 );
and ( n71726 , n71725 , n2667 );
not ( n71727 , n71725 );
and ( n71728 , n71727 , n70007 );
or ( n71729 , n71726 , n71728 );
buf ( n5591 , n71729 );
buf ( n5592 , 1'b0 );
not ( n71732 , n68838 );
buf ( n5594 , n71732 );
buf ( n5595 , n68634 );
and ( n71735 , n71725 , n2623 );
not ( n71736 , n71725 );
and ( n71737 , n71736 , n69947 );
or ( n71738 , n71735 , n71737 );
buf ( n71739 , n71738 );
buf ( n5601 , 1'b0 );
not ( n71741 , n68838 );
buf ( n71742 , n71741 );
buf ( n5604 , n68634 );
and ( n71744 , n71725 , n68770 );
not ( n71745 , n71725 );
not ( n71746 , n69627 );
not ( n71747 , n71746 );
nand ( n71748 , n69896 , n69871 );
nor ( n71749 , n71748 , n69793 );
nand ( n71750 , n71029 , n71749 );
not ( n71751 , n71750 );
not ( n71752 , n69932 );
not ( n71753 , n69850 );
nor ( n71754 , n71752 , n71753 );
not ( n71755 , n71754 );
not ( n71756 , n69685 );
nor ( n71757 , n71755 , n71756 );
nand ( n71758 , n71747 , n71751 , n71757 );
not ( n71759 , n69706 );
and ( n71760 , n71758 , n71759 );
not ( n71761 , n71758 );
and ( n71762 , n71761 , n69706 );
nor ( n71763 , n71760 , n71762 );
and ( n71764 , n71745 , n71763 );
or ( n71765 , n71744 , n71764 );
buf ( n71766 , n71765 );
buf ( n71767 , 1'b0 );
not ( n71768 , n68838 );
buf ( n71769 , n71768 );
buf ( n5631 , n68634 );
and ( n71771 , n71725 , n2633 );
not ( n71772 , n71725 );
not ( n71773 , n71755 );
nand ( n71774 , n71773 , n71751 , n69627 );
and ( n71775 , n71774 , n71756 );
not ( n71776 , n71774 );
and ( n71777 , n71776 , n69685 );
nor ( n71778 , n71775 , n71777 );
not ( n71779 , n71778 );
not ( n71780 , n71779 );
and ( n71781 , n71772 , n71780 );
or ( n71782 , n71771 , n71781 );
buf ( n5644 , n71782 );
buf ( n5645 , 1'b0 );
not ( n71785 , n68838 );
buf ( n71786 , n71785 );
buf ( n71787 , n68634 );
and ( n71788 , n71725 , n2635 );
not ( n71789 , n71725 );
not ( n71790 , n69627 );
not ( n71791 , n71790 );
nand ( n71792 , n71791 , n71751 , n69932 );
and ( n71793 , n71792 , n71753 );
not ( n71794 , n71792 );
not ( n71795 , n71753 );
and ( n71796 , n71794 , n71795 );
nor ( n71797 , n71793 , n71796 );
not ( n71798 , n71797 );
not ( n71799 , n71798 );
and ( n71800 , n71789 , n71799 );
or ( n71801 , n71788 , n71800 );
buf ( n71802 , n71801 );
buf ( n5664 , 1'b0 );
not ( n71804 , n68838 );
buf ( n71805 , n71804 );
buf ( n71806 , n68634 );
and ( n71807 , n71725 , n2637 );
not ( n71808 , n71725 );
nand ( n71809 , n71751 , n69627 );
not ( n71810 , n69932 );
and ( n71811 , n71809 , n71810 );
not ( n71812 , n71809 );
and ( n71813 , n71812 , n69932 );
nor ( n71814 , n71811 , n71813 );
and ( n71815 , n71808 , n71814 );
or ( n71816 , n71807 , n71815 );
buf ( n71817 , n71816 );
buf ( n71818 , 1'b0 );
not ( n71819 , n68838 );
buf ( n5681 , n71819 );
buf ( n5682 , n68634 );
and ( n71822 , n71725 , n2639 );
not ( n71823 , n71725 );
not ( n71824 , n71748 );
nand ( n71825 , n71824 , n69792 );
nor ( n71826 , n71030 , n71825 );
nand ( n71827 , n69627 , n71826 );
not ( n71828 , n69769 );
and ( n71829 , n71827 , n71828 );
not ( n71830 , n71827 );
and ( n71831 , n71830 , n69769 );
nor ( n71832 , n71829 , n71831 );
not ( n71833 , n71832 );
not ( n71834 , n71833 );
and ( n71835 , n71823 , n71834 );
or ( n71836 , n71822 , n71835 );
buf ( n71837 , n71836 );
buf ( n71838 , 1'b0 );
not ( n71839 , n68838 );
buf ( n5701 , n71839 );
buf ( n5702 , n68634 );
not ( n71842 , n71725 );
not ( n71843 , n71842 );
and ( n71844 , n71843 , n68780 );
not ( n71845 , n71843 );
nor ( n71846 , n71030 , n71748 );
nand ( n71847 , n69627 , n71846 );
not ( n71848 , n69792 );
and ( n71849 , n71847 , n71848 );
not ( n71850 , n71847 );
and ( n71851 , n71850 , n69792 );
nor ( n71852 , n71849 , n71851 );
and ( n71853 , n71845 , n71852 );
or ( n71854 , n71844 , n71853 );
buf ( n71855 , n71854 );
buf ( n71856 , 1'b0 );
not ( n71857 , n68838 );
buf ( n71858 , n71857 );
buf ( n71859 , n68634 );
and ( n71860 , n71725 , n2643 );
not ( n71861 , n71725 );
not ( n71862 , n69896 );
and ( n71863 , n71029 , n69871 );
nand ( n71864 , n71863 , n69627 );
not ( n71865 , n71864 );
or ( n71866 , n71862 , n71865 );
nand ( n71867 , n69627 , n71863 );
or ( n71868 , n71867 , n69896 );
nand ( n71869 , n71866 , n71868 );
and ( n71870 , n71861 , n71869 );
or ( n71871 , n71860 , n71870 );
buf ( n71872 , n71871 );
buf ( n5734 , 1'b0 );
not ( n71874 , n68838 );
buf ( n71875 , n71874 );
buf ( n71876 , n68634 );
and ( n71877 , n71843 , n68784 );
not ( n71878 , n71843 );
and ( n71879 , n71878 , n71037 );
or ( n71880 , n71877 , n71879 );
buf ( n5742 , n71880 );
buf ( n71882 , 1'b0 );
not ( n71883 , n68838 );
buf ( n5745 , n71883 );
buf ( n71885 , n68634 );
and ( n71886 , n71843 , n68786 );
not ( n71887 , n71843 );
and ( n71888 , n71887 , n71058 );
or ( n71889 , n71886 , n71888 );
buf ( n5751 , n71889 );
buf ( n5752 , 1'b0 );
not ( n71892 , n68838 );
buf ( n5754 , n71892 );
buf ( n5755 , n68634 );
and ( n71895 , n71843 , n2649 );
not ( n71896 , n71843 );
and ( n71897 , n71896 , n71047 );
or ( n71898 , n71895 , n71897 );
buf ( n71899 , n71898 );
buf ( n71900 , 1'b0 );
not ( n71901 , n68838 );
buf ( n71902 , n71901 );
buf ( n71903 , n68634 );
and ( n71904 , n71843 , n2651 );
not ( n71905 , n71843 );
and ( n71906 , n71905 , n69660 );
or ( n71907 , n71904 , n71906 );
buf ( n71908 , n71907 );
buf ( n71909 , 1'b0 );
not ( n71910 , n68838 );
buf ( n71911 , n71910 );
buf ( n71912 , n68634 );
and ( n71913 , n71843 , n2653 );
not ( n71914 , n71843 );
and ( n71915 , n71914 , n69977 );
or ( n71916 , n71913 , n71915 );
buf ( n71917 , n71916 );
buf ( n71918 , 1'b0 );
not ( n71919 , n68838 );
buf ( n71920 , n71919 );
buf ( n71921 , n68634 );
and ( n71922 , n71725 , n68794 );
not ( n71923 , n71725 );
and ( n71924 , n71923 , n69620 );
or ( n71925 , n71922 , n71924 );
buf ( n71926 , n71925 );
buf ( n71927 , 1'b0 );
not ( n71928 , n68838 );
buf ( n71929 , n71928 );
buf ( n71930 , n68634 );
and ( n71931 , n71725 , n68796 );
not ( n71932 , n71725 );
and ( n71933 , n71932 , n69981 );
or ( n71934 , n71931 , n71933 );
buf ( n71935 , n71934 );
buf ( n71936 , 1'b0 );
not ( n71937 , n68838 );
buf ( n71938 , n71937 );
buf ( n71939 , n68634 );
and ( n71940 , n71725 , n2659 );
not ( n71941 , n71725 );
and ( n71942 , n71941 , n70098 );
or ( n71943 , n71940 , n71942 );
buf ( n71944 , n71943 );
buf ( n71945 , 1'b0 );
not ( n71946 , n68838 );
buf ( n71947 , n71946 );
buf ( n71948 , n68634 );
and ( n71949 , n71725 , n68800 );
not ( n71950 , n71725 );
and ( n71951 , n71950 , n69990 );
or ( n71952 , n71949 , n71951 );
buf ( n71953 , n71952 );
buf ( n71954 , 1'b0 );
not ( n71955 , n68838 );
buf ( n71956 , n71955 );
buf ( n71957 , n68634 );
and ( n71958 , n71725 , n2663 );
not ( n71959 , n71725 );
and ( n71960 , n71959 , n71530 );
or ( n71961 , n71958 , n71960 );
buf ( n71962 , n71961 );
buf ( n71963 , 1'b0 );
not ( n71964 , n68838 );
buf ( n71965 , n71964 );
buf ( n71966 , n68634 );
and ( n71967 , n71725 , n2665 );
not ( n71968 , n71725 );
and ( n71969 , n71968 , n70013 );
or ( n71970 , n71967 , n71969 );
buf ( n71971 , n71970 );
buf ( n71972 , 1'b0 );
not ( n71973 , n68838 );
buf ( n71974 , n71973 );
buf ( n71975 , n68634 );
buf ( n71976 , n70859 );
buf ( n71977 , 1'b0 );
not ( n71978 , n68838 );
buf ( n71979 , n71978 );
buf ( n71980 , n68634 );
not ( n71981 , n70922 );
nand ( n71982 , n70164 , n70180 , n70863 );
and ( n71983 , n70207 , n70139 );
nand ( n71984 , n70136 , n70196 , n71983 );
nor ( n71985 , n71982 , n71984 );
not ( n71986 , n71985 );
or ( n71987 , n71981 , n71986 );
not ( n71988 , n70862 );
nor ( n71989 , n71988 , n71982 );
nand ( n71990 , n71989 , n70571 );
nand ( n71991 , n71989 , n70566 );
not ( n71992 , n70139 );
nor ( n71993 , n71985 , n71992 );
nand ( n71994 , n71990 , n71991 , n71993 );
not ( n71995 , n71994 );
not ( n71996 , n70847 );
not ( n71997 , n71989 );
or ( n71998 , n71996 , n71997 );
nand ( n71999 , n71998 , n70875 );
nand ( n72000 , n70136 , n70872 , n71983 );
nor ( n72001 , n71982 , n72000 );
nor ( n72002 , n71999 , n72001 );
nand ( n72003 , n71995 , n72002 );
not ( n72004 , n72003 );
and ( n72005 , n70883 , n69537 );
not ( n72006 , n70883 );
and ( n72007 , n72006 , n70884 );
nor ( n72008 , n72005 , n72007 );
not ( n72009 , n72008 );
and ( n72010 , n72004 , n72009 );
not ( n72011 , n71991 );
and ( n72012 , n70965 , n72011 );
nor ( n72013 , n72010 , n72012 );
not ( n72014 , n71990 );
and ( n72015 , n70992 , n72014 );
not ( n72016 , n72001 );
not ( n72017 , n72016 );
nand ( n72018 , n71008 , n72017 );
nand ( n72019 , n71999 , n70263 );
nand ( n72020 , n69537 , n70859 );
nand ( n72021 , n72018 , n72019 , n72020 );
nor ( n72022 , n72015 , n72021 );
and ( n72023 , n72013 , n72022 );
nand ( n72024 , n71987 , n72023 );
buf ( n72025 , n72024 );
buf ( n72026 , 1'b0 );
not ( n72027 , n68838 );
buf ( n5889 , n72027 );
buf ( n72029 , n68634 );
not ( n72030 , n69358 );
not ( n72031 , n70007 );
nand ( n72032 , n69971 , n70092 );
not ( n72033 , n72032 );
or ( n72034 , n72031 , n72033 );
or ( n72035 , n72032 , n70007 );
nand ( n72036 , n72034 , n72035 );
not ( n72037 , n72036 );
or ( n72038 , n72030 , n72037 );
nand ( n72039 , n70090 , n71272 );
nand ( n72040 , n72038 , n72039 );
not ( n72041 , n72040 );
or ( n72042 , n72041 , n71986 );
nand ( n72043 , n70641 , n70987 );
not ( n72044 , n72043 );
not ( n72045 , n70984 );
or ( n72046 , n72044 , n72045 );
or ( n72047 , n70984 , n72043 );
nand ( n72048 , n72046 , n72047 );
nand ( n72049 , n72048 , n72014 );
nand ( n72050 , n70392 , n70960 );
not ( n72051 , n72050 );
not ( n72052 , n70957 );
or ( n72053 , n72051 , n72052 );
or ( n72054 , n70957 , n72050 );
nand ( n72055 , n72053 , n72054 );
nand ( n72056 , n72055 , n72011 );
not ( n72057 , n72003 );
and ( n72058 , n70882 , n69549 );
not ( n72059 , n70882 );
not ( n72060 , n69549 );
and ( n72061 , n72059 , n72060 );
nor ( n72062 , n72058 , n72061 );
nand ( n72063 , n72057 , n72062 );
nand ( n72064 , n71999 , n70378 );
not ( n72065 , n70378 );
not ( n72066 , n71003 );
or ( n72067 , n72065 , n72066 );
or ( n72068 , n71003 , n70378 );
nand ( n72069 , n72067 , n72068 );
nand ( n72070 , n72069 , n72017 );
not ( n72071 , n70859 );
nor ( n72072 , n72060 , n72071 );
not ( n72073 , n72072 );
and ( n72074 , n72064 , n72070 , n72073 );
and ( n72075 , n72049 , n72056 , n72063 , n72074 );
nand ( n72076 , n72042 , n72075 );
buf ( n72077 , n72076 );
buf ( n72078 , 1'b0 );
not ( n72079 , n68838 );
buf ( n72080 , n72079 );
buf ( n72081 , n68634 );
and ( n72082 , n71272 , n70031 );
not ( n72083 , n71272 );
not ( n72084 , n70082 );
not ( n72085 , n72084 );
nand ( n72086 , n69971 , n70076 );
not ( n72087 , n70090 );
nor ( n72088 , n72086 , n72087 );
not ( n72089 , n72088 );
or ( n72090 , n72085 , n72089 );
or ( n72091 , n72088 , n72084 );
nand ( n72092 , n72090 , n72091 );
and ( n72093 , n72083 , n72092 );
nor ( n72094 , n72082 , n72093 );
or ( n72095 , n72094 , n71986 );
not ( n72096 , n70480 );
nand ( n72097 , n72096 , n70541 );
not ( n72098 , n72097 );
not ( n72099 , n70495 );
nor ( n72100 , n70936 , n72099 );
not ( n72101 , n72100 );
not ( n72102 , n70947 );
or ( n72103 , n72101 , n72102 );
not ( n72104 , n70950 );
or ( n72105 , n72104 , n72099 );
nand ( n72106 , n72105 , n70488 );
not ( n72107 , n72106 );
nand ( n72108 , n72103 , n72107 );
not ( n72109 , n72108 );
or ( n72110 , n72098 , n72109 );
or ( n72111 , n72108 , n72097 );
nand ( n72112 , n72110 , n72111 );
nand ( n72113 , n72112 , n72011 );
nand ( n72114 , n70617 , n70611 );
not ( n72115 , n72114 );
not ( n72116 , n70616 );
nor ( n72117 , n72116 , n70971 );
not ( n72118 , n72117 );
not ( n72119 , n70978 );
or ( n72120 , n72118 , n72119 );
not ( n72121 , n70616 );
not ( n72122 , n70769 );
or ( n72123 , n72121 , n72122 );
nand ( n72124 , n72123 , n70597 );
not ( n72125 , n72124 );
nand ( n72126 , n72120 , n72125 );
not ( n72127 , n72126 );
or ( n72128 , n72115 , n72127 );
or ( n72129 , n72126 , n72114 );
nand ( n72130 , n72128 , n72129 );
nand ( n72131 , n72130 , n72014 );
and ( n72132 , n70880 , n70881 );
not ( n72133 , n70880 );
and ( n72134 , n72133 , n3324 );
nor ( n72135 , n72132 , n72134 );
nand ( n72136 , n72057 , n72135 );
and ( n72137 , n71999 , n70388 );
nor ( n72138 , n70881 , n72071 );
not ( n72139 , n72138 );
not ( n72140 , n70388 );
not ( n72141 , n71000 );
not ( n72142 , n70432 );
not ( n72143 , n70818 );
nand ( n72144 , n72142 , n72143 );
or ( n72145 , n72144 , n70477 );
nor ( n72146 , n72141 , n72145 );
not ( n72147 , n72146 );
or ( n72148 , n72140 , n72147 );
or ( n72149 , n72146 , n70388 );
nand ( n72150 , n72148 , n72149 );
nand ( n72151 , n72150 , n72017 );
nand ( n72152 , n72139 , n72151 );
nor ( n72153 , n72137 , n72152 );
and ( n72154 , n72113 , n72131 , n72136 , n72153 );
nand ( n72155 , n72095 , n72154 );
buf ( n6017 , n72155 );
buf ( n72157 , 1'b0 );
not ( n72158 , n68838 );
buf ( n72159 , n72158 );
buf ( n6021 , n68634 );
and ( n72161 , n69359 , n70024 );
not ( n72162 , n69359 );
not ( n72163 , n70090 );
not ( n72164 , n72086 );
or ( n72165 , n72163 , n72164 );
or ( n72166 , n72086 , n70090 );
nand ( n72167 , n72165 , n72166 );
and ( n72168 , n72162 , n72167 );
nor ( n72169 , n72161 , n72168 );
or ( n72170 , n72169 , n71986 );
nand ( n72171 , n70616 , n70597 );
not ( n72172 , n72171 );
not ( n72173 , n70769 );
nand ( n72174 , n72173 , n70762 );
not ( n72175 , n72174 );
or ( n72176 , n72172 , n72175 );
or ( n72177 , n72174 , n72171 );
nand ( n72178 , n72176 , n72177 );
nand ( n72179 , n72178 , n72014 );
not ( n72180 , n72099 );
nand ( n72181 , n72180 , n70488 );
not ( n72182 , n72181 );
nor ( n72183 , n70936 , n70462 );
not ( n72184 , n72183 );
not ( n72185 , n70530 );
or ( n72186 , n72184 , n72185 );
nand ( n72187 , n72186 , n72104 );
not ( n72188 , n72187 );
or ( n72189 , n72182 , n72188 );
or ( n72190 , n72187 , n72181 );
nand ( n72191 , n72189 , n72190 );
nand ( n72192 , n72191 , n72011 );
and ( n72193 , n70879 , n3288 );
not ( n72194 , n70879 );
not ( n72195 , n3288 );
and ( n72196 , n72194 , n72195 );
nor ( n72197 , n72193 , n72196 );
nand ( n72198 , n72057 , n72197 );
and ( n72199 , n71999 , n70477 );
nor ( n72200 , n72195 , n72071 );
not ( n72201 , n72200 );
not ( n72202 , n70477 );
nor ( n72203 , n72141 , n72144 );
not ( n72204 , n72203 );
or ( n72205 , n72202 , n72204 );
or ( n72206 , n72203 , n70477 );
nand ( n72207 , n72205 , n72206 );
nand ( n72208 , n72207 , n72017 );
nand ( n72209 , n72201 , n72208 );
nor ( n72210 , n72199 , n72209 );
and ( n72211 , n72179 , n72192 , n72198 , n72210 );
nand ( n72212 , n72170 , n72211 );
buf ( n72213 , n72212 );
buf ( n72214 , 1'b0 );
not ( n72215 , n68838 );
buf ( n6077 , n72215 );
buf ( n72217 , n68634 );
and ( n72218 , n71272 , n70038 );
not ( n72219 , n71272 );
not ( n72220 , n70031 );
not ( n72221 , n70075 );
nand ( n72222 , n72221 , n69971 );
not ( n72223 , n72222 );
nand ( n72224 , n72223 , n70024 );
not ( n72225 , n72224 );
or ( n72226 , n72220 , n72225 );
or ( n72227 , n72224 , n70031 );
nand ( n72228 , n72226 , n72227 );
and ( n72229 , n72219 , n72228 );
nor ( n72230 , n72218 , n72229 );
or ( n72231 , n72230 , n71986 );
nand ( n72232 , n70539 , n70542 );
not ( n72233 , n72232 );
not ( n72234 , n70426 );
not ( n72235 , n72234 );
not ( n72236 , n70947 );
or ( n72237 , n72235 , n72236 );
nand ( n72238 , n72237 , n70535 );
not ( n72239 , n72238 );
or ( n72240 , n72233 , n72239 );
or ( n72241 , n72238 , n72232 );
nand ( n72242 , n72240 , n72241 );
nand ( n72243 , n72242 , n72011 );
nand ( n72244 , n70745 , n70768 );
not ( n72245 , n72244 );
not ( n72246 , n70759 );
not ( n72247 , n70978 );
or ( n72248 , n72246 , n72247 );
not ( n72249 , n70763 );
nand ( n72250 , n72248 , n72249 );
not ( n72251 , n72250 );
or ( n72252 , n72245 , n72251 );
or ( n72253 , n72250 , n72244 );
nand ( n72254 , n72252 , n72253 );
nand ( n72255 , n72254 , n72014 );
and ( n72256 , n70878 , n70877 );
not ( n72257 , n70878 );
and ( n72258 , n72257 , n3356 );
nor ( n72259 , n72256 , n72258 );
nand ( n72260 , n72057 , n72259 );
and ( n72261 , n71999 , n70432 );
nor ( n72262 , n70877 , n72071 );
not ( n72263 , n72262 );
not ( n72264 , n70432 );
nor ( n72265 , n72141 , n70818 );
not ( n72266 , n72265 );
or ( n72267 , n72264 , n72266 );
or ( n72268 , n72265 , n70432 );
nand ( n72269 , n72267 , n72268 );
nand ( n72270 , n72269 , n72017 );
nand ( n72271 , n72263 , n72270 );
nor ( n72272 , n72261 , n72271 );
and ( n72273 , n72243 , n72255 , n72260 , n72272 );
nand ( n72274 , n72231 , n72273 );
buf ( n6136 , n72274 );
buf ( n6137 , 1'b0 );
not ( n72277 , n68838 );
buf ( n72278 , n72277 );
buf ( n72279 , n68634 );
not ( n72280 , n69358 );
not ( n72281 , n70024 );
not ( n72282 , n72222 );
or ( n72283 , n72281 , n72282 );
or ( n72284 , n72222 , n70024 );
nand ( n72285 , n72283 , n72284 );
not ( n72286 , n72285 );
or ( n72287 , n72280 , n72286 );
nand ( n72288 , n70040 , n71272 );
nand ( n72289 , n72287 , n72288 );
not ( n72290 , n72289 );
or ( n72291 , n72290 , n71986 );
nand ( n72292 , n72234 , n70535 );
xnor ( n72293 , n70947 , n72292 );
nand ( n72294 , n72293 , n72011 );
nand ( n72295 , n70759 , n72249 );
not ( n72296 , n72295 );
not ( n72297 , n70978 );
or ( n72298 , n72296 , n72297 );
or ( n72299 , n70978 , n72295 );
nand ( n72300 , n72298 , n72299 );
nand ( n72301 , n72300 , n72014 );
not ( n72302 , n70817 );
and ( n72303 , n71999 , n72302 );
and ( n72304 , n71000 , n72143 );
not ( n72305 , n71000 );
and ( n72306 , n72305 , n70818 );
nor ( n72307 , n72304 , n72306 );
not ( n72308 , n72307 );
not ( n72309 , n72017 );
or ( n72310 , n72308 , n72309 );
nand ( n72311 , n3344 , n70859 );
nand ( n72312 , n72310 , n72311 );
nor ( n72313 , n72303 , n72312 );
nand ( n72314 , n72294 , n72301 , n72313 );
not ( n72315 , n3344 );
and ( n72316 , n72315 , n3304 );
not ( n72317 , n3304 );
and ( n72318 , n72317 , n3344 );
nor ( n72319 , n72316 , n72318 );
nor ( n72320 , n72003 , n72319 );
nor ( n72321 , n72314 , n72320 );
nand ( n72322 , n72291 , n72321 );
buf ( n6184 , n72322 );
buf ( n6185 , 1'b0 );
not ( n72325 , n68838 );
buf ( n72326 , n72325 );
buf ( n72327 , n68634 );
and ( n72328 , n69359 , n70073 );
not ( n72329 , n69359 );
not ( n72330 , n70073 );
nand ( n72331 , n69969 , n70053 );
nor ( n72332 , n72330 , n72331 );
nand ( n72333 , n72332 , n70040 );
not ( n72334 , n70038 );
and ( n72335 , n72333 , n72334 );
not ( n72336 , n72333 );
and ( n72337 , n72336 , n70038 );
nor ( n72338 , n72335 , n72337 );
and ( n72339 , n72329 , n72338 );
nor ( n72340 , n72328 , n72339 );
or ( n72341 , n72340 , n71986 );
not ( n72342 , n70940 );
nand ( n72343 , n72342 , n70528 );
nand ( n72344 , n70463 , n70527 );
xnor ( n72345 , n72343 , n72344 );
and ( n72346 , n72345 , n72011 );
and ( n72347 , n71999 , n70420 );
nor ( n72348 , n72346 , n72347 );
not ( n72349 , n70974 );
nand ( n72350 , n72349 , n70733 );
not ( n72351 , n72350 );
nand ( n72352 , n70761 , n70732 );
not ( n72353 , n72352 );
or ( n72354 , n72351 , n72353 );
or ( n72355 , n72352 , n72350 );
nand ( n72356 , n72354 , n72355 );
and ( n72357 , n72356 , n72014 );
not ( n72358 , n72017 );
not ( n72359 , n70420 );
not ( n72360 , n70831 );
nor ( n72361 , n72360 , n70459 );
not ( n72362 , n72361 );
or ( n72363 , n72359 , n72362 );
or ( n72364 , n72361 , n70420 );
nand ( n72365 , n72363 , n72364 );
not ( n72366 , n72365 );
or ( n72367 , n72358 , n72366 );
nor ( n72368 , n72317 , n72071 );
not ( n72369 , n72368 );
nand ( n72370 , n72367 , n72369 );
nor ( n72371 , n72357 , n72370 );
nand ( n72372 , n72057 , n72317 );
and ( n72373 , n72348 , n72371 , n72372 );
nand ( n72374 , n72341 , n72373 );
buf ( n72375 , n72374 );
buf ( n72376 , 1'b0 );
not ( n72377 , n68838 );
buf ( n72378 , n72377 );
buf ( n72379 , n68634 );
and ( n72380 , n71272 , n70053 );
not ( n72381 , n71272 );
xor ( n72382 , n70040 , n72332 );
and ( n72383 , n72381 , n72382 );
nor ( n72384 , n72380 , n72383 );
or ( n72385 , n72384 , n71986 );
nand ( n72386 , n72003 , n72071 );
and ( n72387 , n72386 , n3915 );
not ( n72388 , n72016 );
not ( n72389 , n70459 );
not ( n72390 , n70831 );
or ( n72391 , n72389 , n72390 );
or ( n72392 , n70831 , n70459 );
nand ( n72393 , n72391 , n72392 );
not ( n72394 , n72393 );
not ( n72395 , n72394 );
and ( n72396 , n72388 , n72395 );
not ( n72397 , n70516 );
nand ( n72398 , n72397 , n70528 );
not ( n72399 , n72398 );
or ( n72400 , n70507 , n70524 );
nand ( n72401 , n72400 , n70518 );
not ( n72402 , n72401 );
or ( n72403 , n72399 , n72402 );
or ( n72404 , n72398 , n72401 );
nand ( n72405 , n72403 , n72404 );
and ( n72406 , n72405 , n72011 );
nor ( n72407 , n72396 , n72406 );
not ( n72408 , n71999 );
not ( n72409 , n72408 );
not ( n72410 , n70459 );
not ( n72411 , n72410 );
and ( n72412 , n72409 , n72411 );
not ( n72413 , n70727 );
nand ( n72414 , n70716 , n70733 );
not ( n72415 , n72414 );
or ( n72416 , n72413 , n72415 );
or ( n72417 , n72414 , n70727 );
nand ( n72418 , n72416 , n72417 );
and ( n72419 , n72418 , n72014 );
nor ( n72420 , n72412 , n72419 );
nand ( n72421 , n72407 , n72420 );
nor ( n72422 , n72387 , n72421 );
nand ( n72423 , n72385 , n72422 );
buf ( n72424 , n72423 );
buf ( n72425 , 1'b0 );
not ( n72426 , n68838 );
buf ( n72427 , n72426 );
buf ( n72428 , n68634 );
and ( n72429 , n71272 , n71763 );
not ( n72430 , n71272 );
not ( n72431 , n71814 );
nand ( n72432 , n71852 , n71832 );
nor ( n72433 , n72431 , n72432 );
and ( n72434 , n71587 , n72433 , n71520 );
nand ( n72435 , n71037 , n71869 );
not ( n72436 , n72435 );
nand ( n72437 , n69660 , n71058 );
not ( n72438 , n72437 );
nand ( n72439 , n69977 , n70098 );
nor ( n72440 , n69982 , n72439 );
nand ( n72441 , n72436 , n72438 , n72440 , n71047 );
nor ( n72442 , n69970 , n72441 );
not ( n72443 , n71763 );
nand ( n72444 , n71797 , n71778 );
nor ( n72445 , n72443 , n72444 );
nand ( n72446 , n72434 , n72442 , n72445 );
not ( n72447 , n71746 );
not ( n72448 , n69707 );
nand ( n72449 , n72448 , n71754 );
not ( n72450 , n72449 );
nand ( n72451 , n72447 , n71751 , n72450 );
xnor ( n72452 , n72451 , n69729 );
not ( n72453 , n72452 );
nor ( n72454 , n72446 , n72453 );
not ( n72455 , n72454 );
not ( n72456 , n69743 );
not ( n72457 , n69729 );
nor ( n72458 , n72457 , n72449 );
nand ( n72459 , n72447 , n71751 , n72458 );
not ( n72460 , n72459 );
or ( n72461 , n72456 , n72460 );
or ( n72462 , n72459 , n69743 );
nand ( n72463 , n72461 , n72462 );
not ( n72464 , n72463 );
and ( n72465 , n72455 , n72464 );
not ( n72466 , n72455 );
and ( n72467 , n72466 , n72463 );
nor ( n72468 , n72465 , n72467 );
and ( n72469 , n72430 , n72468 );
nor ( n72470 , n72429 , n72469 );
or ( n72471 , n72470 , n71986 );
nor ( n72472 , n71131 , n71100 );
and ( n72473 , n72472 , n71085 );
nand ( n72474 , n70222 , n68646 );
not ( n72475 , n72474 );
not ( n72476 , n72475 );
not ( n72477 , n72476 );
not ( n72478 , n69896 );
not ( n72479 , n72478 );
or ( n72480 , n72477 , n72479 );
nand ( n72481 , n69896 , n72475 );
nand ( n72482 , n72480 , n72481 );
not ( n72483 , n69871 );
nand ( n72484 , n70222 , n2508 );
not ( n72485 , n72484 );
nor ( n72486 , n72483 , n72485 );
nor ( n72487 , n72482 , n72486 );
not ( n72488 , n72485 );
not ( n72489 , n69871 );
or ( n72490 , n72488 , n72489 );
not ( n72491 , n72485 );
not ( n72492 , n69871 );
nand ( n72493 , n72491 , n72492 );
nand ( n72494 , n72490 , n72493 );
nor ( n72495 , n71126 , n71122 );
nor ( n72496 , n72494 , n72495 );
nor ( n72497 , n72487 , n72496 );
nand ( n72498 , n70222 , n68645 );
not ( n72499 , n72498 );
not ( n72500 , n72499 );
not ( n72501 , n69792 );
or ( n72502 , n72500 , n72501 );
not ( n72503 , n72499 );
not ( n72504 , n69792 );
nand ( n72505 , n72503 , n72504 );
nand ( n72506 , n72502 , n72505 );
and ( n72507 , n69896 , n72476 );
nor ( n72508 , n72506 , n72507 );
nand ( n72509 , n70222 , n68644 );
not ( n72510 , n72509 );
not ( n72511 , n72510 );
not ( n72512 , n69769 );
or ( n72513 , n72511 , n72512 );
not ( n72514 , n69769 );
not ( n72515 , n72510 );
nand ( n72516 , n72514 , n72515 );
nand ( n72517 , n72513 , n72516 );
nor ( n72518 , n72504 , n72499 );
nor ( n72519 , n72517 , n72518 );
nor ( n72520 , n72508 , n72519 );
and ( n72521 , n72497 , n72520 );
nand ( n72522 , n72473 , n72521 );
and ( n72523 , n70222 , n2501 );
not ( n72524 , n72523 );
not ( n72525 , n69706 );
or ( n72526 , n72524 , n72525 );
not ( n72527 , n72523 );
not ( n72528 , n69706 );
nand ( n72529 , n72527 , n72528 );
nand ( n72530 , n72526 , n72529 );
not ( n72531 , n69685 );
not ( n72532 , n71070 );
nand ( n72533 , n72532 , n2502 );
not ( n72534 , n72533 );
nor ( n72535 , n72531 , n72534 );
nor ( n72536 , n72530 , n72535 );
not ( n72537 , n72534 );
not ( n72538 , n69685 );
or ( n72539 , n72537 , n72538 );
not ( n72540 , n72534 );
not ( n72541 , n69685 );
nand ( n72542 , n72540 , n72541 );
nand ( n72543 , n72539 , n72542 );
and ( n72544 , n70222 , n2503 );
not ( n72545 , n72544 );
and ( n72546 , n69850 , n72545 );
nor ( n72547 , n72543 , n72546 );
nor ( n72548 , n72536 , n72547 );
not ( n72549 , n72544 );
not ( n72550 , n69850 );
or ( n72551 , n72549 , n72550 );
not ( n72552 , n69850 );
nand ( n72553 , n72552 , n72545 );
nand ( n72554 , n72551 , n72553 );
not ( n72555 , n69932 );
nand ( n72556 , n72532 , n2504 );
not ( n72557 , n72556 );
nor ( n72558 , n72555 , n72557 );
nor ( n72559 , n72554 , n72558 );
not ( n72560 , n72557 );
not ( n72561 , n69932 );
or ( n72562 , n72560 , n72561 );
not ( n72563 , n72557 );
not ( n72564 , n69932 );
nand ( n72565 , n72563 , n72564 );
nand ( n72566 , n72562 , n72565 );
and ( n72567 , n69769 , n72515 );
nor ( n72568 , n72566 , n72567 );
nor ( n72569 , n72559 , n72568 );
nand ( n72570 , n72548 , n72569 );
nor ( n72571 , n72522 , n72570 );
not ( n72572 , n72571 );
not ( n72573 , n70553 );
or ( n72574 , n72572 , n72573 );
not ( n72575 , n72570 );
not ( n72576 , n72575 );
not ( n72577 , n72521 );
not ( n72578 , n71109 );
not ( n72579 , n72472 );
or ( n72580 , n72578 , n72579 );
not ( n72581 , n71131 );
not ( n72582 , n71112 );
and ( n72583 , n72581 , n72582 );
nor ( n72584 , n72583 , n71132 );
nand ( n72585 , n72580 , n72584 );
not ( n72586 , n72585 );
or ( n72587 , n72577 , n72586 );
not ( n72588 , n72520 );
and ( n72589 , n72494 , n72495 );
not ( n72590 , n72589 );
not ( n72591 , n72487 );
not ( n72592 , n72591 );
or ( n72593 , n72590 , n72592 );
nand ( n72594 , n72482 , n72486 );
nand ( n72595 , n72593 , n72594 );
not ( n72596 , n72595 );
or ( n72597 , n72588 , n72596 );
nand ( n72598 , n72506 , n72507 );
nor ( n72599 , n72519 , n72598 );
and ( n72600 , n72517 , n72518 );
nor ( n72601 , n72599 , n72600 );
nand ( n72602 , n72597 , n72601 );
not ( n72603 , n72602 );
nand ( n72604 , n72587 , n72603 );
not ( n72605 , n72604 );
or ( n72606 , n72576 , n72605 );
not ( n72607 , n72548 );
nand ( n72608 , n72566 , n72567 );
or ( n72609 , n72559 , n72608 );
nand ( n72610 , n72554 , n72558 );
nand ( n72611 , n72609 , n72610 );
not ( n72612 , n72611 );
or ( n72613 , n72607 , n72612 );
not ( n72614 , n72536 );
nand ( n72615 , n72543 , n72546 );
not ( n72616 , n72615 );
and ( n72617 , n72614 , n72616 );
and ( n72618 , n72530 , n72535 );
nor ( n72619 , n72617 , n72618 );
nand ( n72620 , n72613 , n72619 );
not ( n72621 , n72620 );
nand ( n72622 , n72606 , n72621 );
not ( n72623 , n72622 );
nand ( n72624 , n72574 , n72623 );
nand ( n72625 , n70222 , n2500 );
not ( n72626 , n72625 );
not ( n72627 , n72626 );
not ( n72628 , n69729 );
not ( n72629 , n72628 );
not ( n72630 , n72629 );
or ( n72631 , n72627 , n72630 );
not ( n72632 , n72626 );
not ( n72633 , n72629 );
nand ( n72634 , n72632 , n72633 );
nand ( n72635 , n72631 , n72634 );
not ( n72636 , n69706 );
nor ( n72637 , n72636 , n72523 );
nor ( n72638 , n72635 , n72637 );
not ( n72639 , n72638 );
nand ( n72640 , n72635 , n72637 );
nand ( n72641 , n72639 , n72640 );
not ( n72642 , n72641 );
and ( n72643 , n72624 , n72642 );
not ( n72644 , n72624 );
and ( n72645 , n72644 , n72641 );
nor ( n72646 , n72643 , n72645 );
nand ( n72647 , n72646 , n72011 );
xor ( n72648 , n72523 , n69706 );
and ( n72649 , n69685 , n72534 );
nor ( n72650 , n72648 , n72649 );
not ( n72651 , n69685 );
not ( n72652 , n72534 );
not ( n72653 , n72652 );
or ( n72654 , n72651 , n72653 );
not ( n72655 , n69685 );
nand ( n72656 , n72655 , n72534 );
nand ( n72657 , n72654 , n72656 );
and ( n72658 , n72544 , n69850 );
nor ( n72659 , n72657 , n72658 );
nor ( n72660 , n72650 , n72659 );
xor ( n72661 , n72544 , n69850 );
and ( n72662 , n69932 , n72557 );
nor ( n72663 , n72661 , n72662 );
not ( n72664 , n72557 );
not ( n72665 , n72664 );
not ( n72666 , n69932 );
or ( n72667 , n72665 , n72666 );
not ( n72668 , n69932 );
nand ( n72669 , n72668 , n72557 );
nand ( n72670 , n72667 , n72669 );
and ( n72671 , n69769 , n72510 );
nor ( n72672 , n72670 , n72671 );
nor ( n72673 , n72663 , n72672 );
and ( n72674 , n72660 , n72673 );
not ( n72675 , n72674 );
not ( n72676 , n72475 );
not ( n72677 , n69896 );
not ( n72678 , n72677 );
or ( n72679 , n72676 , n72678 );
not ( n72680 , n72475 );
nand ( n72681 , n72680 , n69896 );
nand ( n72682 , n72679 , n72681 );
and ( n72683 , n69871 , n72485 );
nor ( n72684 , n72682 , n72683 );
not ( n72685 , n72684 );
not ( n72686 , n72485 );
not ( n72687 , n69871 );
not ( n72688 , n72687 );
or ( n72689 , n72686 , n72688 );
not ( n72690 , n72485 );
nand ( n72691 , n72690 , n69871 );
nand ( n72692 , n72689 , n72691 );
not ( n72693 , n72692 );
and ( n72694 , n69804 , n71122 );
not ( n72695 , n72694 );
nand ( n72696 , n72693 , n72695 );
nand ( n72697 , n72685 , n72696 );
not ( n72698 , n72697 );
not ( n72699 , n72499 );
not ( n72700 , n69792 );
not ( n72701 , n72700 );
or ( n72702 , n72699 , n72701 );
not ( n72703 , n72499 );
nand ( n72704 , n69792 , n72703 );
nand ( n72705 , n72702 , n72704 );
and ( n72706 , n69896 , n72475 );
nor ( n72707 , n72705 , n72706 );
not ( n72708 , n72510 );
not ( n72709 , n72708 );
not ( n72710 , n69769 );
or ( n72711 , n72709 , n72710 );
not ( n72712 , n69769 );
nand ( n72713 , n72712 , n72510 );
nand ( n72714 , n72711 , n72713 );
nand ( n72715 , n69792 , n72499 );
not ( n72716 , n72715 );
nor ( n72717 , n72714 , n72716 );
nor ( n72718 , n72707 , n72717 );
nand ( n72719 , n72698 , n72718 );
not ( n72720 , n72719 );
nor ( n72721 , n71169 , n71146 );
not ( n72722 , n72721 );
nor ( n72723 , n72722 , n71160 );
nand ( n72724 , n72720 , n72723 );
nor ( n72725 , n72675 , n72724 );
not ( n72726 , n72725 );
not ( n72727 , n70809 );
or ( n72728 , n72726 , n72727 );
nand ( n72729 , n72705 , n72706 );
or ( n72730 , n72717 , n72729 );
nand ( n72731 , n72714 , n72716 );
nand ( n72732 , n72730 , n72731 );
not ( n72733 , n72732 );
not ( n72734 , n72718 );
and ( n72735 , n72733 , n72734 );
nand ( n72736 , n72692 , n72694 );
or ( n72737 , n72684 , n72736 );
nand ( n72738 , n72682 , n72683 );
nand ( n72739 , n72737 , n72738 );
nor ( n72740 , n72732 , n72739 );
and ( n72741 , n72740 , n72697 );
nor ( n72742 , n72735 , n72741 );
nand ( n72743 , n71178 , n72721 );
not ( n72744 , n71146 );
not ( n72745 , n71181 );
and ( n72746 , n72744 , n72745 );
nor ( n72747 , n72746 , n71145 );
nand ( n72748 , n72740 , n72743 , n72747 );
nand ( n72749 , n72742 , n72748 );
not ( n72750 , n72749 );
and ( n72751 , n72750 , n72674 );
not ( n72752 , n72660 );
nand ( n72753 , n72670 , n72671 );
or ( n72754 , n72663 , n72753 );
nand ( n72755 , n72661 , n72662 );
nand ( n72756 , n72754 , n72755 );
not ( n72757 , n72756 );
or ( n72758 , n72752 , n72757 );
not ( n72759 , n72650 );
nand ( n72760 , n72657 , n72658 );
not ( n72761 , n72760 );
and ( n72762 , n72759 , n72761 );
nand ( n72763 , n72648 , n72649 );
not ( n72764 , n72763 );
nor ( n72765 , n72762 , n72764 );
nand ( n72766 , n72758 , n72765 );
nor ( n72767 , n72751 , n72766 );
nand ( n72768 , n72728 , n72767 );
xor ( n72769 , n72626 , n69729 );
and ( n72770 , n72523 , n69706 );
or ( n72771 , n72769 , n72770 );
nand ( n72772 , n72769 , n72770 );
nand ( n72773 , n72771 , n72772 );
not ( n72774 , n72773 );
and ( n72775 , n72768 , n72774 );
not ( n72776 , n72768 );
and ( n72777 , n72776 , n72773 );
nor ( n72778 , n72775 , n72777 );
and ( n72779 , n72778 , n72014 );
not ( n72780 , n69720 );
not ( n72781 , n69702 );
nor ( n72782 , n70893 , n70894 );
nand ( n72783 , n72782 , n3514 );
not ( n72784 , n69818 );
nor ( n72785 , n72783 , n72784 );
nand ( n72786 , n72785 , n69802 );
not ( n72787 , n69851 );
nor ( n72788 , n72786 , n72787 );
and ( n72789 , n72788 , n69887 );
nand ( n72790 , n72789 , n69772 );
not ( n72791 , n69766 );
nor ( n72792 , n72790 , n72791 );
nand ( n72793 , n72792 , n69928 );
not ( n72794 , n3707 );
nor ( n72795 , n72793 , n72794 );
nand ( n72796 , n72795 , n69676 );
nor ( n72797 , n72781 , n72796 );
not ( n72798 , n72797 );
or ( n72799 , n72780 , n72798 );
or ( n72800 , n72797 , n69720 );
nand ( n72801 , n72799 , n72800 );
not ( n72802 , n72801 );
or ( n72803 , n72802 , n72003 );
not ( n72804 , n72626 );
not ( n72805 , n71092 );
not ( n72806 , n71122 );
nand ( n72807 , n72805 , n72806 );
nor ( n72808 , n72807 , n71194 );
nor ( n72809 , n72499 , n72510 );
nor ( n72810 , n72485 , n72475 );
and ( n72811 , n72809 , n72810 );
and ( n72812 , n72808 , n72811 );
nor ( n72813 , n72557 , n72544 );
not ( n72814 , n72523 );
not ( n72815 , n72814 );
nor ( n72816 , n72815 , n72534 );
and ( n72817 , n72813 , n72816 );
nand ( n72818 , n72812 , n72817 );
nor ( n72819 , n70832 , n72818 );
not ( n72820 , n72819 );
or ( n72821 , n72804 , n72820 );
or ( n72822 , n72819 , n72626 );
nand ( n72823 , n72821 , n72822 );
nand ( n72824 , n72823 , n72017 );
nand ( n72825 , n71999 , n72626 );
nand ( n72826 , n69721 , n70859 );
and ( n72827 , n72824 , n72825 , n72826 );
nand ( n72828 , n72803 , n72827 );
nor ( n72829 , n72779 , n72828 );
and ( n72830 , n72647 , n72829 );
nand ( n72831 , n72471 , n72830 );
buf ( n72832 , n72831 );
buf ( n72833 , 1'b0 );
not ( n72834 , n68838 );
buf ( n6696 , n72834 );
buf ( n72836 , n68634 );
and ( n72837 , n69359 , n71780 );
not ( n72838 , n69359 );
and ( n72839 , n72446 , n72453 );
not ( n72840 , n72446 );
not ( n72841 , n72453 );
and ( n72842 , n72840 , n72841 );
nor ( n72843 , n72839 , n72842 );
and ( n72844 , n72838 , n72843 );
nor ( n72845 , n72837 , n72844 );
or ( n72846 , n72845 , n71986 );
not ( n72847 , n72547 );
and ( n72848 , n72569 , n72847 );
not ( n72849 , n72848 );
nor ( n72850 , n72522 , n72849 );
not ( n72851 , n72850 );
not ( n72852 , n70553 );
or ( n72853 , n72851 , n72852 );
not ( n72854 , n72848 );
not ( n72855 , n72604 );
or ( n72856 , n72854 , n72855 );
not ( n72857 , n72847 );
not ( n72858 , n72611 );
or ( n72859 , n72857 , n72858 );
nand ( n72860 , n72859 , n72615 );
not ( n72861 , n72860 );
nand ( n72862 , n72856 , n72861 );
not ( n72863 , n72862 );
nand ( n72864 , n72853 , n72863 );
or ( n72865 , n72536 , n72618 );
xnor ( n72866 , n72864 , n72865 );
nand ( n72867 , n72866 , n72011 );
not ( n72868 , n72650 );
nand ( n72869 , n72868 , n72763 );
not ( n72870 , n72869 );
not ( n72871 , n72659 );
nand ( n72872 , n72673 , n72871 );
nor ( n72873 , n72724 , n72872 );
not ( n72874 , n72873 );
not ( n72875 , n70804 );
or ( n72876 , n72874 , n72875 );
not ( n72877 , n72749 );
not ( n72878 , n72872 );
and ( n72879 , n72877 , n72878 );
not ( n72880 , n72871 );
not ( n72881 , n72756 );
or ( n72882 , n72880 , n72881 );
nand ( n72883 , n72882 , n72760 );
nor ( n72884 , n72879 , n72883 );
nand ( n72885 , n72876 , n72884 );
not ( n72886 , n72885 );
or ( n72887 , n72870 , n72886 );
or ( n72888 , n72885 , n72869 );
nand ( n72889 , n72887 , n72888 );
and ( n72890 , n72889 , n72014 );
and ( n72891 , n72796 , n69702 );
not ( n72892 , n72796 );
and ( n72893 , n72892 , n69701 );
nor ( n72894 , n72891 , n72893 );
or ( n72895 , n72003 , n72894 );
not ( n72896 , n72815 );
not ( n72897 , n72557 );
nor ( n72898 , n72807 , n70225 );
nor ( n72899 , n72544 , n72534 );
and ( n72900 , n72809 , n72899 , n71193 );
nand ( n72901 , n72897 , n72898 , n72900 , n72810 );
nor ( n72902 , n70832 , n72901 );
not ( n72903 , n72902 );
or ( n72904 , n72896 , n72903 );
or ( n72905 , n72902 , n72815 );
nand ( n72906 , n72904 , n72905 );
and ( n72907 , n72906 , n72017 );
nor ( n72908 , n69701 , n72071 );
nor ( n72909 , n72907 , n72908 );
nand ( n72910 , n71999 , n72815 );
nand ( n72911 , n72895 , n72909 , n72910 );
nor ( n72912 , n72890 , n72911 );
and ( n72913 , n72867 , n72912 );
nand ( n72914 , n72846 , n72913 );
buf ( n6776 , n72914 );
buf ( n6777 , 1'b0 );
not ( n72917 , n68838 );
buf ( n72918 , n72917 );
buf ( n72919 , n68634 );
and ( n72920 , n71272 , n71799 );
not ( n72921 , n71272 );
not ( n72922 , n72441 );
nand ( n72923 , n72922 , n72434 );
not ( n72924 , n72923 );
not ( n72925 , n72444 );
nand ( n72926 , n72924 , n69969 , n72925 );
not ( n72927 , n71763 );
and ( n72928 , n72926 , n72927 );
not ( n72929 , n72926 );
and ( n72930 , n72929 , n71763 );
nor ( n72931 , n72928 , n72930 );
and ( n72932 , n72921 , n72931 );
nor ( n72933 , n72920 , n72932 );
or ( n72934 , n72933 , n71986 );
not ( n72935 , n72569 );
nor ( n72936 , n72935 , n72522 );
not ( n72937 , n72936 );
not ( n72938 , n70553 );
or ( n72939 , n72937 , n72938 );
not ( n72940 , n72569 );
not ( n72941 , n72604 );
or ( n72942 , n72940 , n72941 );
not ( n72943 , n72611 );
nand ( n72944 , n72942 , n72943 );
not ( n72945 , n72944 );
nand ( n72946 , n72939 , n72945 );
nand ( n72947 , n72847 , n72615 );
not ( n72948 , n72947 );
and ( n72949 , n72946 , n72948 );
not ( n72950 , n72946 );
and ( n72951 , n72950 , n72947 );
nor ( n72952 , n72949 , n72951 );
nand ( n72953 , n72952 , n72011 );
not ( n72954 , n72673 );
nor ( n72955 , n72724 , n72954 );
not ( n72956 , n72955 );
not ( n72957 , n70804 );
or ( n72958 , n72956 , n72957 );
and ( n72959 , n72750 , n72673 );
nor ( n72960 , n72959 , n72756 );
nand ( n72961 , n72958 , n72960 );
nand ( n72962 , n72871 , n72760 );
not ( n72963 , n72962 );
and ( n72964 , n72961 , n72963 );
not ( n72965 , n72961 );
and ( n72966 , n72965 , n72962 );
nor ( n72967 , n72964 , n72966 );
and ( n72968 , n72967 , n72014 );
and ( n72969 , n72795 , n69675 );
not ( n72970 , n72795 );
and ( n72971 , n72970 , n69676 );
nor ( n72972 , n72969 , n72971 );
or ( n72973 , n72003 , n72972 );
not ( n72974 , n72534 );
not ( n72975 , n72807 );
not ( n72976 , n71194 );
nand ( n72977 , n72975 , n72976 , n72811 , n72813 );
nor ( n72978 , n70832 , n72977 );
not ( n72979 , n72978 );
or ( n72980 , n72974 , n72979 );
or ( n72981 , n72978 , n72534 );
nand ( n72982 , n72980 , n72981 );
and ( n72983 , n72982 , n72017 );
nor ( n72984 , n69675 , n72071 );
nor ( n72985 , n72983 , n72984 );
nand ( n72986 , n71999 , n72534 );
nand ( n72987 , n72973 , n72985 , n72986 );
nor ( n72988 , n72968 , n72987 );
and ( n72989 , n72953 , n72988 );
nand ( n72990 , n72934 , n72989 );
buf ( n6852 , n72990 );
buf ( n72992 , 1'b0 );
not ( n72993 , n68838 );
buf ( n72994 , n72993 );
buf ( n6856 , n68634 );
and ( n72996 , n69359 , n71814 );
not ( n72997 , n69359 );
not ( n72998 , n69969 );
nor ( n72999 , n72923 , n72998 );
nand ( n73000 , n72999 , n71797 );
not ( n73001 , n71778 );
and ( n73002 , n73000 , n73001 );
not ( n73003 , n73000 );
and ( n73004 , n73003 , n71778 );
nor ( n73005 , n73002 , n73004 );
and ( n73006 , n72997 , n73005 );
nor ( n73007 , n72996 , n73006 );
or ( n73008 , n73007 , n71986 );
nor ( n73009 , n72522 , n72568 );
not ( n73010 , n73009 );
not ( n73011 , n70553 );
or ( n73012 , n73010 , n73011 );
not ( n73013 , n72568 );
not ( n73014 , n73013 );
not ( n73015 , n72604 );
or ( n73016 , n73014 , n73015 );
nand ( n73017 , n73016 , n72608 );
not ( n73018 , n73017 );
nand ( n73019 , n73012 , n73018 );
not ( n73020 , n72559 );
nand ( n73021 , n73020 , n72610 );
xnor ( n73022 , n73019 , n73021 );
nand ( n73023 , n73022 , n72011 );
not ( n73024 , n72663 );
nand ( n73025 , n73024 , n72755 );
not ( n73026 , n73025 );
nor ( n73027 , n72724 , n72672 );
not ( n73028 , n73027 );
not ( n73029 , n70804 );
or ( n73030 , n73028 , n73029 );
not ( n73031 , n72749 );
not ( n73032 , n72672 );
and ( n73033 , n73031 , n73032 );
not ( n73034 , n72753 );
nor ( n73035 , n73033 , n73034 );
nand ( n73036 , n73030 , n73035 );
not ( n73037 , n73036 );
or ( n73038 , n73026 , n73037 );
or ( n73039 , n73036 , n73025 );
nand ( n73040 , n73038 , n73039 );
and ( n73041 , n73040 , n72014 );
and ( n73042 , n72793 , n3707 );
not ( n73043 , n72793 );
and ( n73044 , n73043 , n72794 );
nor ( n73045 , n73042 , n73044 );
or ( n73046 , n72003 , n73045 );
not ( n73047 , n72544 );
not ( n73048 , n72499 );
and ( n73049 , n72810 , n73048 );
nor ( n73050 , n71074 , n72557 , n72510 );
nand ( n73051 , n72898 , n73049 , n73050 );
nor ( n73052 , n70832 , n73051 );
not ( n73053 , n73052 );
or ( n73054 , n73047 , n73053 );
or ( n73055 , n73052 , n72544 );
nand ( n73056 , n73054 , n73055 );
and ( n73057 , n73056 , n72017 );
nor ( n73058 , n72794 , n72071 );
nor ( n73059 , n73057 , n73058 );
nand ( n73060 , n71999 , n72544 );
nand ( n73061 , n73046 , n73059 , n73060 );
nor ( n73062 , n73041 , n73061 );
and ( n73063 , n73023 , n73062 );
nand ( n73064 , n73008 , n73063 );
buf ( n6926 , n73064 );
buf ( n6927 , 1'b0 );
not ( n73067 , n68838 );
buf ( n73068 , n73067 );
buf ( n73069 , n68634 );
and ( n73070 , n71272 , n71834 );
not ( n73071 , n71272 );
not ( n73072 , n72999 );
not ( n73073 , n71797 );
and ( n73074 , n73072 , n73073 );
not ( n73075 , n73072 );
and ( n73076 , n73075 , n71797 );
nor ( n73077 , n73074 , n73076 );
and ( n73078 , n73071 , n73077 );
nor ( n73079 , n73070 , n73078 );
or ( n73080 , n73079 , n71986 );
not ( n73081 , n72522 );
not ( n73082 , n73081 );
not ( n73083 , n70553 );
or ( n73084 , n73082 , n73083 );
not ( n73085 , n72604 );
nand ( n73086 , n73084 , n73085 );
nand ( n73087 , n73013 , n72608 );
not ( n73088 , n73087 );
and ( n73089 , n73086 , n73088 );
not ( n73090 , n73086 );
and ( n73091 , n73090 , n73087 );
nor ( n73092 , n73089 , n73091 );
nand ( n73093 , n73092 , n72011 );
not ( n73094 , n72724 );
not ( n73095 , n73094 );
not ( n73096 , n70809 );
or ( n73097 , n73095 , n73096 );
nand ( n73098 , n73097 , n72749 );
nor ( n73099 , n73034 , n72672 );
and ( n73100 , n73098 , n73099 );
not ( n73101 , n73098 );
not ( n73102 , n73099 );
and ( n73103 , n73101 , n73102 );
nor ( n73104 , n73100 , n73103 );
and ( n73105 , n73104 , n72014 );
and ( n73106 , n72792 , n69927 );
not ( n73107 , n72792 );
and ( n73108 , n73107 , n69928 );
nor ( n73109 , n73106 , n73108 );
or ( n73110 , n72003 , n73109 );
not ( n73111 , n72557 );
not ( n73112 , n72812 );
nor ( n73113 , n73112 , n70832 );
not ( n73114 , n73113 );
or ( n73115 , n73111 , n73114 );
or ( n73116 , n73113 , n72557 );
nand ( n73117 , n73115 , n73116 );
and ( n73118 , n73117 , n72017 );
nor ( n73119 , n69927 , n72071 );
nor ( n73120 , n73118 , n73119 );
nand ( n73121 , n71999 , n72557 );
nand ( n73122 , n73110 , n73120 , n73121 );
nor ( n73123 , n73105 , n73122 );
and ( n73124 , n73093 , n73123 );
nand ( n73125 , n73080 , n73124 );
buf ( n6987 , n73125 );
buf ( n73127 , 1'b0 );
not ( n73128 , n68838 );
buf ( n73129 , n73128 );
buf ( n6991 , n68634 );
and ( n73131 , n69359 , n71852 );
not ( n73132 , n69359 );
nor ( n73133 , n72441 , n71522 );
nand ( n73134 , n73133 , n71852 );
not ( n73135 , n73134 );
nand ( n73136 , n73135 , n71832 );
not ( n73137 , n71814 );
and ( n73138 , n73136 , n73137 );
not ( n73139 , n73136 );
and ( n73140 , n73139 , n71814 );
nor ( n73141 , n73138 , n73140 );
and ( n73142 , n73132 , n73141 );
nor ( n73143 , n73131 , n73142 );
or ( n73144 , n73143 , n71986 );
not ( n73145 , n72473 );
not ( n73146 , n72508 );
and ( n73147 , n72497 , n73146 );
not ( n73148 , n73147 );
nor ( n73149 , n73145 , n73148 );
not ( n73150 , n73149 );
not ( n73151 , n70553 );
or ( n73152 , n73150 , n73151 );
and ( n73153 , n73147 , n72585 );
not ( n73154 , n73146 );
not ( n73155 , n72595 );
or ( n73156 , n73154 , n73155 );
nand ( n73157 , n73156 , n72598 );
nor ( n73158 , n73153 , n73157 );
nand ( n73159 , n73152 , n73158 );
or ( n73160 , n72600 , n72519 );
xnor ( n73161 , n73159 , n73160 );
nand ( n73162 , n73161 , n72011 );
not ( n73163 , n72717 );
nand ( n73164 , n73163 , n72731 );
not ( n73165 , n73164 );
nor ( n73166 , n72697 , n72707 );
not ( n73167 , n73166 );
not ( n73168 , n72723 );
nor ( n73169 , n73167 , n73168 );
not ( n73170 , n73169 );
not ( n73171 , n70809 );
or ( n73172 , n73170 , n73171 );
not ( n73173 , n73166 );
nand ( n73174 , n72743 , n72747 );
not ( n73175 , n73174 );
or ( n73176 , n73173 , n73175 );
not ( n73177 , n72707 );
not ( n73178 , n73177 );
not ( n73179 , n72739 );
or ( n73180 , n73178 , n73179 );
nand ( n73181 , n73180 , n72729 );
not ( n73182 , n73181 );
nand ( n73183 , n73176 , n73182 );
not ( n73184 , n73183 );
nand ( n73185 , n73172 , n73184 );
not ( n73186 , n73185 );
or ( n73187 , n73165 , n73186 );
or ( n73188 , n73185 , n73164 );
nand ( n73189 , n73187 , n73188 );
and ( n73190 , n73189 , n72014 );
and ( n73191 , n72790 , n69766 );
not ( n73192 , n72790 );
and ( n73193 , n73192 , n72791 );
nor ( n73194 , n73191 , n73193 );
or ( n73195 , n72003 , n73194 );
not ( n73196 , n72510 );
nand ( n73197 , n72808 , n73049 );
nor ( n73198 , n70832 , n73197 );
not ( n73199 , n73198 );
or ( n73200 , n73196 , n73199 );
or ( n73201 , n73198 , n72510 );
nand ( n73202 , n73200 , n73201 );
and ( n73203 , n73202 , n72017 );
nor ( n73204 , n72791 , n72071 );
nor ( n73205 , n73203 , n73204 );
nand ( n73206 , n71999 , n72510 );
nand ( n73207 , n73195 , n73205 , n73206 );
nor ( n73208 , n73190 , n73207 );
and ( n73209 , n73162 , n73208 );
nand ( n73210 , n73144 , n73209 );
buf ( n73211 , n73210 );
buf ( n73212 , 1'b0 );
not ( n73213 , n68838 );
buf ( n73214 , n73213 );
buf ( n73215 , n68634 );
and ( n73216 , n71272 , n71869 );
not ( n73217 , n71272 );
not ( n73218 , n71832 );
and ( n73219 , n73134 , n73218 );
not ( n73220 , n73134 );
and ( n73221 , n73220 , n71832 );
nor ( n73222 , n73219 , n73221 );
and ( n73223 , n73217 , n73222 );
nor ( n73224 , n73216 , n73223 );
or ( n73225 , n73224 , n71986 );
not ( n73226 , n72497 );
nor ( n73227 , n73145 , n73226 );
not ( n73228 , n73227 );
not ( n73229 , n70553 );
or ( n73230 , n73228 , n73229 );
and ( n73231 , n72497 , n72585 );
nor ( n73232 , n73231 , n72595 );
nand ( n73233 , n73230 , n73232 );
nand ( n73234 , n73146 , n72598 );
not ( n73235 , n73234 );
and ( n73236 , n73233 , n73235 );
not ( n73237 , n73233 );
and ( n73238 , n73237 , n73234 );
nor ( n73239 , n73236 , n73238 );
nand ( n73240 , n73239 , n72011 );
nor ( n73241 , n73168 , n72697 );
not ( n73242 , n73241 );
not ( n73243 , n70809 );
or ( n73244 , n73242 , n73243 );
and ( n73245 , n72698 , n73174 );
nor ( n73246 , n73245 , n72739 );
nand ( n73247 , n73244 , n73246 );
nand ( n73248 , n73177 , n72729 );
not ( n73249 , n73248 );
and ( n73250 , n73247 , n73249 );
not ( n73251 , n73247 );
and ( n73252 , n73251 , n73248 );
nor ( n73253 , n73250 , n73252 );
and ( n73254 , n73253 , n72014 );
and ( n73255 , n72789 , n69771 );
not ( n73256 , n72789 );
and ( n73257 , n73256 , n69772 );
nor ( n73258 , n73255 , n73257 );
or ( n73259 , n72003 , n73258 );
not ( n73260 , n72499 );
nand ( n73261 , n72808 , n72810 );
nor ( n73262 , n70832 , n73261 );
not ( n73263 , n73262 );
or ( n73264 , n73260 , n73263 );
or ( n73265 , n73262 , n72499 );
nand ( n73266 , n73264 , n73265 );
and ( n73267 , n73266 , n72017 );
nor ( n73268 , n69771 , n72071 );
nor ( n73269 , n73267 , n73268 );
nand ( n73270 , n71999 , n72499 );
nand ( n73271 , n73259 , n73269 , n73270 );
nor ( n73272 , n73254 , n73271 );
and ( n73273 , n73240 , n73272 );
nand ( n73274 , n73225 , n73273 );
buf ( n73275 , n73274 );
buf ( n73276 , 1'b0 );
not ( n73277 , n68838 );
buf ( n7139 , n73277 );
buf ( n73279 , n68634 );
and ( n73280 , n69359 , n71037 );
not ( n73281 , n69359 );
not ( n73282 , n71852 );
not ( n73283 , n73133 );
not ( n73284 , n73283 );
or ( n73285 , n73282 , n73284 );
or ( n73286 , n71852 , n73283 );
nand ( n73287 , n73285 , n73286 );
and ( n73288 , n73281 , n73287 );
nor ( n73289 , n73280 , n73288 );
or ( n73290 , n73289 , n71986 );
nor ( n73291 , n73145 , n72496 );
not ( n73292 , n73291 );
not ( n73293 , n70553 );
or ( n73294 , n73292 , n73293 );
not ( n73295 , n72496 );
not ( n73296 , n73295 );
not ( n73297 , n72585 );
or ( n73298 , n73296 , n73297 );
not ( n73299 , n72589 );
nand ( n73300 , n73298 , n73299 );
not ( n73301 , n73300 );
nand ( n73302 , n73294 , n73301 );
nand ( n73303 , n72591 , n72594 );
xnor ( n73304 , n73302 , n73303 );
nand ( n73305 , n73304 , n72011 );
not ( n73306 , n72684 );
nand ( n73307 , n73306 , n72738 );
not ( n73308 , n73307 );
not ( n73309 , n72696 );
nor ( n73310 , n73309 , n73168 );
not ( n73311 , n73310 );
not ( n73312 , n70809 );
or ( n73313 , n73311 , n73312 );
not ( n73314 , n72696 );
not ( n73315 , n73174 );
or ( n73316 , n73314 , n73315 );
nand ( n73317 , n73316 , n72736 );
not ( n73318 , n73317 );
nand ( n73319 , n73313 , n73318 );
not ( n73320 , n73319 );
or ( n73321 , n73308 , n73320 );
or ( n73322 , n73319 , n73307 );
nand ( n73323 , n73321 , n73322 );
and ( n73324 , n72014 , n73323 );
and ( n73325 , n72788 , n69886 );
not ( n73326 , n72788 );
and ( n73327 , n73326 , n69887 );
nor ( n73328 , n73325 , n73327 );
or ( n73329 , n72003 , n73328 );
not ( n73330 , n72475 );
not ( n73331 , n72485 );
nand ( n73332 , n73331 , n72808 );
nor ( n73333 , n70832 , n73332 );
not ( n73334 , n73333 );
or ( n73335 , n73330 , n73334 );
or ( n73336 , n73333 , n72475 );
nand ( n73337 , n73335 , n73336 );
and ( n73338 , n73337 , n72017 );
nor ( n73339 , n69886 , n72071 );
nor ( n73340 , n73338 , n73339 );
nand ( n73341 , n71999 , n72475 );
nand ( n73342 , n73329 , n73340 , n73341 );
nor ( n73343 , n73324 , n73342 );
and ( n73344 , n73305 , n73343 );
nand ( n73345 , n73290 , n73344 );
buf ( n7207 , n73345 );
buf ( n7208 , 1'b0 );
not ( n73348 , n68838 );
buf ( n73349 , n73348 );
buf ( n73350 , n68634 );
and ( n73351 , n71272 , n71058 );
not ( n73352 , n71272 );
not ( n73353 , n71059 );
nand ( n73354 , n73353 , n71037 );
not ( n73355 , n71869 );
and ( n73356 , n73354 , n73355 );
not ( n73357 , n73354 );
and ( n73358 , n73357 , n71869 );
nor ( n73359 , n73356 , n73358 );
and ( n73360 , n73352 , n73359 );
nor ( n73361 , n73351 , n73360 );
or ( n73362 , n73361 , n71986 );
not ( n73363 , n72473 );
not ( n73364 , n70553 );
or ( n73365 , n73363 , n73364 );
not ( n73366 , n72585 );
nand ( n73367 , n73365 , n73366 );
nand ( n73368 , n73295 , n73299 );
xnor ( n73369 , n73367 , n73368 );
nand ( n73370 , n73369 , n72011 );
nand ( n73371 , n72696 , n72736 );
not ( n73372 , n73371 );
not ( n73373 , n72723 );
not ( n73374 , n70809 );
or ( n73375 , n73373 , n73374 );
not ( n73376 , n73174 );
nand ( n73377 , n73375 , n73376 );
not ( n73378 , n73377 );
or ( n73379 , n73372 , n73378 );
or ( n73380 , n73377 , n73371 );
nand ( n73381 , n73379 , n73380 );
and ( n73382 , n73381 , n72014 );
and ( n73383 , n72786 , n69851 );
not ( n73384 , n72786 );
and ( n73385 , n73384 , n72787 );
nor ( n73386 , n73383 , n73385 );
or ( n73387 , n72003 , n73386 );
not ( n73388 , n72485 );
not ( n73389 , n72808 );
nor ( n73390 , n70832 , n73389 );
not ( n73391 , n73390 );
or ( n73392 , n73388 , n73391 );
or ( n73393 , n73390 , n72485 );
nand ( n73394 , n73392 , n73393 );
and ( n73395 , n73394 , n72017 );
nor ( n73396 , n72787 , n72071 );
nor ( n73397 , n73395 , n73396 );
nand ( n73398 , n71999 , n72485 );
nand ( n73399 , n73387 , n73397 , n73398 );
nor ( n73400 , n73382 , n73399 );
and ( n73401 , n73370 , n73400 );
nand ( n73402 , n73362 , n73401 );
buf ( n73403 , n73402 );
buf ( n73404 , 1'b0 );
not ( n73405 , n68838 );
buf ( n73406 , n73405 );
buf ( n73407 , n68634 );
and ( n73408 , n71272 , n69967 );
not ( n73409 , n71272 );
not ( n73410 , n70073 );
not ( n73411 , n72331 );
or ( n73412 , n73410 , n73411 );
or ( n73413 , n72331 , n70073 );
nand ( n73414 , n73412 , n73413 );
and ( n73415 , n73409 , n73414 );
nor ( n73416 , n73408 , n73415 );
or ( n73417 , n73416 , n71986 );
and ( n73418 , n72386 , n70041 );
not ( n73419 , n70524 );
not ( n73420 , n73419 );
not ( n73421 , n70507 );
nand ( n73422 , n73421 , n70518 );
not ( n73423 , n73422 );
or ( n73424 , n73420 , n73423 );
or ( n73425 , n73422 , n73419 );
nand ( n73426 , n73424 , n73425 );
nand ( n73427 , n73426 , n72011 );
xor ( n73428 , n70722 , n70725 );
nand ( n73429 , n72014 , n73428 );
nand ( n73430 , n71999 , n70503 );
not ( n73431 , n70829 );
not ( n73432 , n70522 );
or ( n73433 , n73431 , n73432 );
or ( n73434 , n70522 , n70829 );
nand ( n73435 , n73433 , n73434 );
nand ( n73436 , n72017 , n73435 );
nand ( n73437 , n73427 , n73429 , n73430 , n73436 );
nor ( n73438 , n73418 , n73437 );
nand ( n73439 , n73417 , n73438 );
buf ( n73440 , n73439 );
buf ( n73441 , 1'b0 );
not ( n73442 , n68838 );
buf ( n73443 , n73442 );
buf ( n7305 , n68634 );
not ( n73445 , n71067 );
or ( n73446 , n73445 , n71986 );
nand ( n73447 , n71134 , n72011 );
and ( n73448 , n71188 , n72014 );
not ( n73449 , n69802 );
and ( n73450 , n72785 , n73449 );
not ( n73451 , n72785 );
and ( n73452 , n73451 , n69802 );
nor ( n73453 , n73450 , n73452 );
or ( n73454 , n72003 , n73453 );
and ( n73455 , n71200 , n72017 );
nor ( n73456 , n73449 , n72071 );
nor ( n73457 , n73455 , n73456 );
nand ( n73458 , n71999 , n71122 );
nand ( n73459 , n73454 , n73457 , n73458 );
nor ( n73460 , n73448 , n73459 );
and ( n73461 , n73447 , n73460 );
nand ( n73462 , n73446 , n73461 );
buf ( n73463 , n73462 );
buf ( n73464 , 1'b0 );
not ( n73465 , n68838 );
buf ( n7327 , n73465 );
buf ( n7328 , n68634 );
not ( n73468 , n71225 );
or ( n73469 , n73468 , n71986 );
nand ( n73470 , n71233 , n72011 );
and ( n73471 , n71248 , n72014 );
and ( n73472 , n72783 , n69818 );
not ( n73473 , n72783 );
and ( n73474 , n73473 , n72784 );
nor ( n73475 , n73472 , n73474 );
or ( n73476 , n72003 , n73475 );
and ( n73477 , n71256 , n72017 );
nor ( n73478 , n72784 , n72071 );
nor ( n73479 , n73477 , n73478 );
nand ( n73480 , n71999 , n71092 );
nand ( n73481 , n73476 , n73479 , n73480 );
nor ( n73482 , n73471 , n73481 );
and ( n73483 , n73470 , n73482 );
nand ( n73484 , n73469 , n73483 );
buf ( n73485 , n73484 );
buf ( n73486 , 1'b0 );
not ( n73487 , n68838 );
buf ( n7349 , n73487 );
buf ( n7350 , n68634 );
or ( n73490 , n71281 , n71986 );
nand ( n73491 , n71291 , n72011 );
and ( n73492 , n71304 , n72014 );
not ( n73493 , n3514 );
and ( n73494 , n72782 , n73493 );
not ( n73495 , n72782 );
and ( n73496 , n73495 , n3514 );
nor ( n73497 , n73494 , n73496 );
or ( n73498 , n72003 , n73497 );
and ( n73499 , n71312 , n72017 );
nor ( n73500 , n73493 , n72071 );
nor ( n73501 , n73499 , n73500 );
nand ( n73502 , n71999 , n71074 );
nand ( n73503 , n73498 , n73501 , n73502 );
nor ( n73504 , n73492 , n73503 );
and ( n73505 , n73491 , n73504 );
nand ( n73506 , n73490 , n73505 );
buf ( n73507 , n73506 );
buf ( n73508 , 1'b0 );
not ( n73509 , n68838 );
buf ( n73510 , n73509 );
buf ( n73511 , n68634 );
or ( n73512 , n70109 , n71986 );
not ( n73513 , n70557 );
not ( n73514 , n73513 );
not ( n73515 , n71991 );
and ( n73516 , n73514 , n73515 );
nand ( n73517 , n70812 , n72014 );
nand ( n73518 , n72057 , n70898 );
nand ( n73519 , n70837 , n72017 );
nand ( n73520 , n71999 , n70225 );
nor ( n73521 , n70894 , n72071 );
not ( n73522 , n73521 );
and ( n73523 , n73519 , n73520 , n73522 );
nand ( n73524 , n73517 , n73518 , n73523 );
nor ( n73525 , n73516 , n73524 );
nand ( n73526 , n73512 , n73525 );
buf ( n7388 , n73526 );
buf ( n7389 , 1'b0 );
not ( n73529 , n68838 );
buf ( n7391 , n73529 );
buf ( n7392 , n68634 );
not ( n73532 , n71364 );
or ( n73533 , n73532 , n71986 );
not ( n73534 , n72003 );
not ( n73535 , n69603 );
and ( n73536 , n70892 , n73535 );
not ( n73537 , n70892 );
and ( n73538 , n73537 , n69603 );
nor ( n73539 , n73536 , n73538 );
not ( n73540 , n73539 );
and ( n73541 , n73534 , n73540 );
and ( n73542 , n71390 , n72011 );
nor ( n73543 , n73541 , n73542 );
and ( n73544 , n72014 , n71416 );
nand ( n73545 , n71428 , n72017 );
nand ( n73546 , n71999 , n70238 );
nand ( n73547 , n69603 , n70859 );
nand ( n73548 , n73545 , n73546 , n73547 );
nor ( n73549 , n73544 , n73548 );
and ( n73550 , n73543 , n73549 );
nand ( n73551 , n73533 , n73550 );
buf ( n73552 , n73551 );
buf ( n73553 , 1'b0 );
not ( n73554 , n68838 );
buf ( n73555 , n73554 );
buf ( n73556 , n68634 );
not ( n73557 , n71457 );
or ( n73558 , n73557 , n71986 );
not ( n73559 , n72003 );
and ( n73560 , n70890 , n3454 );
not ( n73561 , n70890 );
and ( n73562 , n73561 , n70891 );
nor ( n73563 , n73560 , n73562 );
not ( n73564 , n73563 );
and ( n73565 , n73559 , n73564 );
and ( n73566 , n71475 , n72011 );
nor ( n73567 , n73565 , n73566 );
and ( n73568 , n72014 , n71491 );
nand ( n73569 , n71501 , n72017 );
nand ( n73570 , n71999 , n70327 );
nand ( n73571 , n3454 , n70859 );
nand ( n73572 , n73569 , n73570 , n73571 );
nor ( n73573 , n73568 , n73572 );
and ( n73574 , n73567 , n73573 );
nand ( n73575 , n73558 , n73574 );
buf ( n73576 , n73575 );
buf ( n73577 , 1'b0 );
not ( n73578 , n68838 );
buf ( n73579 , n73578 );
buf ( n73580 , n68634 );
not ( n73581 , n69358 );
not ( n73582 , n69981 );
not ( n73583 , n71447 );
or ( n73584 , n73582 , n73583 );
or ( n73585 , n71447 , n69981 );
nand ( n73586 , n73584 , n73585 );
not ( n73587 , n73586 );
or ( n73588 , n73581 , n73587 );
nand ( n73589 , n69990 , n69359 );
nand ( n73590 , n73588 , n73589 );
not ( n73591 , n73590 );
or ( n73592 , n73591 , n71986 );
not ( n73593 , n72003 );
not ( n73594 , n69567 );
and ( n73595 , n70889 , n73594 );
not ( n73596 , n70889 );
and ( n73597 , n73596 , n69567 );
nor ( n73598 , n73595 , n73597 );
not ( n73599 , n73598 );
and ( n73600 , n73593 , n73599 );
nand ( n73601 , n70354 , n70357 );
not ( n73602 , n73601 );
nor ( n73603 , n71372 , n70320 );
not ( n73604 , n73603 );
not ( n73605 , n70957 );
or ( n73606 , n73604 , n73605 );
or ( n73607 , n71377 , n70320 );
nand ( n73608 , n73607 , n70351 );
not ( n73609 , n73608 );
nand ( n73610 , n73606 , n73609 );
not ( n73611 , n73610 );
or ( n73612 , n73602 , n73611 );
or ( n73613 , n73610 , n73601 );
nand ( n73614 , n73612 , n73613 );
and ( n73615 , n73614 , n72011 );
nor ( n73616 , n73600 , n73615 );
not ( n73617 , n70670 );
nand ( n73618 , n73617 , n70786 );
not ( n73619 , n73618 );
nor ( n73620 , n71397 , n70679 );
not ( n73621 , n73620 );
not ( n73622 , n70984 );
or ( n73623 , n73621 , n73622 );
not ( n73624 , n71402 );
not ( n73625 , n70679 );
and ( n73626 , n73624 , n73625 );
not ( n73627 , n70784 );
nor ( n73628 , n73626 , n73627 );
nand ( n73629 , n73623 , n73628 );
not ( n73630 , n73629 );
or ( n73631 , n73619 , n73630 );
or ( n73632 , n73629 , n73618 );
nand ( n73633 , n73631 , n73632 );
and ( n73634 , n72014 , n73633 );
not ( n73635 , n70296 );
not ( n73636 , n73635 );
and ( n73637 , n70827 , n71561 );
nand ( n73638 , n71003 , n73637 );
not ( n73639 , n73638 );
or ( n73640 , n73636 , n73639 );
or ( n73641 , n73638 , n73635 );
nand ( n73642 , n73640 , n73641 );
nand ( n73643 , n73642 , n72017 );
nand ( n73644 , n71999 , n70296 );
nand ( n73645 , n69567 , n70859 );
nand ( n73646 , n73643 , n73644 , n73645 );
nor ( n73647 , n73634 , n73646 );
and ( n73648 , n73616 , n73647 );
nand ( n73649 , n73592 , n73648 );
buf ( n73650 , n73649 );
buf ( n73651 , 1'b0 );
not ( n73652 , n68838 );
buf ( n73653 , n73652 );
buf ( n73654 , n68634 );
not ( n73655 , n71532 );
or ( n73656 , n73655 , n71986 );
not ( n73657 , n72003 );
not ( n73658 , n3442 );
and ( n73659 , n70888 , n73658 );
not ( n73660 , n70888 );
and ( n73661 , n73660 , n3442 );
nor ( n73662 , n73659 , n73661 );
not ( n73663 , n73662 );
and ( n73664 , n73657 , n73663 );
and ( n73665 , n71545 , n72011 );
nor ( n73666 , n73664 , n73665 );
and ( n73667 , n71558 , n72014 );
nand ( n73668 , n71567 , n72017 );
nand ( n73669 , n71999 , n70308 );
nand ( n73670 , n3442 , n70859 );
nand ( n73671 , n73668 , n73669 , n73670 );
nor ( n73672 , n73667 , n73671 );
and ( n73673 , n73666 , n73672 );
nand ( n73674 , n73656 , n73673 );
buf ( n7536 , n73674 );
buf ( n7537 , 1'b0 );
not ( n73677 , n68838 );
buf ( n7539 , n73677 );
buf ( n7540 , n68634 );
not ( n73680 , n71598 );
or ( n73681 , n73680 , n71986 );
not ( n73682 , n72003 );
and ( n73683 , n70886 , n69512 );
not ( n73684 , n70886 );
and ( n73685 , n73684 , n70887 );
nor ( n73686 , n73683 , n73685 );
not ( n73687 , n73686 );
and ( n73688 , n73682 , n73687 );
and ( n73689 , n71618 , n72011 );
nor ( n73690 , n73688 , n73689 );
and ( n73691 , n72014 , n71638 );
nand ( n73692 , n71647 , n72017 );
nand ( n73693 , n71999 , n70273 );
nand ( n73694 , n69512 , n70859 );
nand ( n73695 , n73692 , n73693 , n73694 );
nor ( n73696 , n73691 , n73695 );
and ( n73697 , n73690 , n73696 );
nand ( n73698 , n73681 , n73697 );
buf ( n73699 , n73698 );
buf ( n73700 , 1'b0 );
not ( n73701 , n68838 );
buf ( n73702 , n73701 );
buf ( n73703 , n68634 );
not ( n73704 , n71672 );
or ( n73705 , n73704 , n71986 );
not ( n73706 , n72003 );
not ( n73707 , n69520 );
and ( n73708 , n70885 , n73707 );
not ( n73709 , n70885 );
and ( n73710 , n73709 , n69520 );
nor ( n73711 , n73708 , n73710 );
not ( n73712 , n73711 );
and ( n73713 , n73706 , n73712 );
and ( n73714 , n71685 , n72011 );
nor ( n73715 , n73713 , n73714 );
and ( n73716 , n72014 , n71699 );
nand ( n73717 , n71707 , n72017 );
nand ( n73718 , n71999 , n70253 );
nand ( n73719 , n69520 , n70859 );
nand ( n73720 , n73717 , n73718 , n73719 );
nor ( n73721 , n73716 , n73720 );
and ( n73722 , n73715 , n73721 );
nand ( n73723 , n73705 , n73722 );
buf ( n73724 , n73723 );
buf ( n73725 , 1'b0 );
not ( n73726 , n68838 );
buf ( n73727 , n73726 );
buf ( n73728 , n68634 );
not ( n73729 , n70053 );
not ( n73730 , n69970 );
or ( n73731 , n73729 , n73730 );
not ( n73732 , n70053 );
nand ( n73733 , n73732 , n69971 );
nand ( n73734 , n73731 , n73733 );
nand ( n73735 , n73734 , n69358 );
or ( n73736 , n73735 , n71986 );
nand ( n73737 , n72386 , n69950 );
not ( n73738 , n70522 );
nor ( n73739 , n73738 , n72002 );
not ( n73740 , n70523 );
not ( n73741 , n69967 );
or ( n73742 , n73740 , n73741 );
not ( n73743 , n70523 );
nand ( n73744 , n73743 , n70519 );
nand ( n73745 , n73742 , n73744 );
not ( n73746 , n73745 );
not ( n73747 , n72011 );
or ( n73748 , n73746 , n73747 );
not ( n73749 , n70724 );
not ( n73750 , n69967 );
or ( n73751 , n73749 , n73750 );
or ( n73752 , n69967 , n70724 );
nand ( n73753 , n73751 , n73752 );
nand ( n73754 , n72014 , n73753 );
nand ( n73755 , n73748 , n73754 );
nor ( n73756 , n73739 , n73755 );
nand ( n73757 , n73736 , n73737 , n73756 );
buf ( n7619 , n73757 );
buf ( n73759 , 1'b0 );
not ( n73760 , n68838 );
buf ( n7622 , n73760 );
buf ( n7623 , n68634 );
or ( n73763 , n71981 , n70210 );
and ( n73764 , n70573 , n70992 );
not ( n73765 , n70840 );
not ( n73766 , n73765 );
nand ( n73767 , n71008 , n73766 );
not ( n73768 , n70875 );
not ( n73769 , n72008 );
and ( n73770 , n73768 , n73769 );
and ( n73771 , n70849 , n70263 );
nor ( n73772 , n73770 , n73771 );
nand ( n73773 , n70870 , n69533 );
nand ( n73774 , n73767 , n73772 , n73773 );
nor ( n73775 , n73764 , n73774 );
nand ( n73776 , n70965 , n70568 );
and ( n73777 , n73775 , n73776 );
nand ( n73778 , n73763 , n73777 );
buf ( n7640 , n73778 );
buf ( n7641 , 1'b0 );
not ( n73781 , n68838 );
buf ( n73782 , n73781 );
buf ( n73783 , n68634 );
or ( n73784 , n72041 , n70210 );
nand ( n73785 , n72048 , n70573 );
nand ( n73786 , n72055 , n70568 );
not ( n73787 , n72069 );
not ( n73788 , n70840 );
or ( n73789 , n73787 , n73788 );
and ( n73790 , n70870 , n3405 );
and ( n73791 , n70876 , n72062 );
nor ( n73792 , n73790 , n73791 );
nand ( n73793 , n73789 , n73792 );
not ( n73794 , n70378 );
nor ( n73795 , n70848 , n73794 );
nor ( n73796 , n73793 , n73795 );
and ( n73797 , n73785 , n73786 , n73796 );
nand ( n73798 , n73784 , n73797 );
buf ( n73799 , n73798 );
buf ( n73800 , 1'b0 );
not ( n73801 , n68838 );
buf ( n73802 , n73801 );
buf ( n73803 , n68634 );
or ( n73804 , n72094 , n70210 );
nand ( n73805 , n72112 , n70568 );
nand ( n73806 , n72130 , n70573 );
and ( n73807 , n70849 , n70388 );
and ( n73808 , n70876 , n72135 );
nor ( n73809 , n73807 , n73808 );
nand ( n73810 , n70840 , n72150 );
nand ( n73811 , n70870 , n3320 );
and ( n73812 , n73809 , n73810 , n73811 );
and ( n73813 , n73805 , n73806 , n73812 );
nand ( n73814 , n73804 , n73813 );
buf ( n7676 , n73814 );
buf ( n7677 , 1'b0 );
not ( n73817 , n68838 );
buf ( n73818 , n73817 );
buf ( n73819 , n68634 );
or ( n73820 , n72169 , n70210 );
nand ( n73821 , n72178 , n70573 );
nand ( n73822 , n72191 , n70568 );
and ( n73823 , n70849 , n70477 );
and ( n73824 , n70876 , n72197 );
nor ( n73825 , n73823 , n73824 );
nand ( n73826 , n70840 , n72207 );
nand ( n73827 , n70870 , n3276 );
and ( n73828 , n73825 , n73826 , n73827 );
and ( n73829 , n73821 , n73822 , n73828 );
nand ( n73830 , n73820 , n73829 );
buf ( n7692 , n73830 );
buf ( n7693 , 1'b0 );
not ( n73833 , n68838 );
buf ( n73834 , n73833 );
buf ( n7696 , n68634 );
or ( n73836 , n72230 , n70210 );
nand ( n73837 , n72242 , n70568 );
nand ( n73838 , n72254 , n70573 );
and ( n73839 , n70849 , n70432 );
and ( n73840 , n70876 , n72259 );
nor ( n73841 , n73839 , n73840 );
nand ( n73842 , n70840 , n72269 );
not ( n73843 , n70870 );
not ( n73844 , n73843 );
nand ( n73845 , n73844 , n3350 );
and ( n73846 , n73841 , n73842 , n73845 );
and ( n73847 , n73837 , n73838 , n73846 );
nand ( n73848 , n73836 , n73847 );
buf ( n73849 , n73848 );
buf ( n73850 , 1'b0 );
not ( n73851 , n68838 );
buf ( n73852 , n73851 );
buf ( n7714 , n68634 );
or ( n73854 , n72290 , n70210 );
and ( n73855 , n72300 , n70573 );
not ( n73856 , n3346 );
nor ( n73857 , n73843 , n73856 );
nor ( n73858 , n73855 , n73857 );
nand ( n73859 , n72293 , n70568 );
not ( n73860 , n72302 );
not ( n73861 , n70849 );
or ( n73862 , n73860 , n73861 );
not ( n73863 , n70876 );
or ( n73864 , n73863 , n72319 );
nand ( n73865 , n73862 , n73864 );
not ( n73866 , n70840 );
not ( n73867 , n72307 );
nor ( n73868 , n73866 , n73867 );
nor ( n73869 , n73865 , n73868 );
and ( n73870 , n73858 , n73859 , n73869 );
nand ( n73871 , n73854 , n73870 );
buf ( n73872 , n73871 );
buf ( n73873 , 1'b0 );
not ( n73874 , n68838 );
buf ( n73875 , n73874 );
buf ( n73876 , n68634 );
or ( n73877 , n72340 , n70210 );
nand ( n73878 , n72345 , n70568 );
nand ( n73879 , n72356 , n70573 );
nand ( n73880 , n73766 , n72365 );
and ( n73881 , n70849 , n70420 );
and ( n73882 , n70876 , n72317 );
nor ( n73883 , n73881 , n73882 );
nand ( n73884 , n70870 , n69437 );
and ( n73885 , n73880 , n73883 , n73884 );
and ( n73886 , n73878 , n73879 , n73885 );
nand ( n73887 , n73877 , n73886 );
buf ( n7749 , n73887 );
buf ( n7750 , 1'b0 );
not ( n73890 , n68838 );
buf ( n73891 , n73890 );
buf ( n73892 , n68634 );
and ( n73893 , n70870 , n69940 );
not ( n73894 , n70870 );
not ( n73895 , n69947 );
nand ( n73896 , n72454 , n72463 );
not ( n73897 , n73896 );
not ( n73898 , n71750 );
nor ( n73899 , n72449 , n69744 );
nand ( n73900 , n73898 , n72447 , n73899 );
not ( n73901 , n69908 );
xor ( n73902 , n73900 , n73901 );
nand ( n73903 , n73897 , n73902 );
not ( n73904 , n73903 );
or ( n73905 , n73895 , n73904 );
or ( n73906 , n69947 , n73903 );
nand ( n73907 , n73905 , n73906 );
or ( n73908 , n71272 , n70151 );
nand ( n73909 , n73908 , n70222 );
and ( n73910 , n70196 , n73909 );
nand ( n73911 , n73907 , n73910 );
and ( n73912 , n70222 , n68636 );
not ( n73913 , n73912 );
and ( n73914 , n70222 , n2498 );
not ( n73915 , n73914 );
and ( n73916 , n70222 , n2499 );
nor ( n73917 , n72626 , n73916 );
nand ( n73918 , n73915 , n72812 , n73917 , n72817 );
nor ( n73919 , n70832 , n73918 );
not ( n73920 , n73919 );
or ( n73921 , n73913 , n73920 );
or ( n73922 , n73919 , n73912 );
nand ( n73923 , n73921 , n73922 );
and ( n73924 , n73923 , n70995 );
not ( n73925 , n73912 );
nor ( n73926 , n73925 , n70846 );
nor ( n73927 , n73924 , n73926 );
nand ( n73928 , n73911 , n73927 );
and ( n73929 , n73894 , n73928 );
or ( n73930 , n73893 , n73929 );
buf ( n73931 , n73930 );
buf ( n7793 , 1'b0 );
not ( n73933 , n68838 );
buf ( n73934 , n73933 );
buf ( n73935 , n68634 );
and ( n73936 , n70870 , n69902 );
not ( n73937 , n70870 );
and ( n73938 , n70847 , n73914 );
not ( n73939 , n73914 );
nand ( n73940 , n72812 , n72817 , n73917 );
nor ( n73941 , n70832 , n73940 );
not ( n73942 , n73941 );
or ( n73943 , n73939 , n73942 );
or ( n73944 , n73941 , n73914 );
nand ( n73945 , n73943 , n73944 );
and ( n73946 , n73945 , n70995 );
nor ( n73947 , n73938 , n73946 );
nand ( n73948 , n73911 , n73947 );
and ( n73949 , n73937 , n73948 );
or ( n73950 , n73936 , n73949 );
buf ( n73951 , n73950 );
buf ( n73952 , 1'b0 );
not ( n73953 , n68838 );
buf ( n73954 , n73953 );
buf ( n73955 , n68634 );
or ( n73956 , n72384 , n70210 );
nand ( n73957 , n72405 , n70568 );
nand ( n73958 , n70573 , n72418 );
nand ( n73959 , n70876 , n3915 );
nand ( n73960 , n73957 , n73958 , n73959 );
or ( n73961 , n73765 , n72394 );
not ( n73962 , n70058 );
or ( n73963 , n73843 , n73962 );
or ( n73964 , n70848 , n72410 );
nand ( n73965 , n73961 , n73963 , n73964 );
nor ( n73966 , n73960 , n73965 );
nand ( n73967 , n73956 , n73966 );
buf ( n7829 , n73967 );
buf ( n7830 , 1'b0 );
not ( n73970 , n68838 );
buf ( n7832 , n73970 );
buf ( n7833 , n68634 );
not ( n73973 , n73902 );
not ( n73974 , n73973 );
not ( n73975 , n73897 );
or ( n73976 , n73974 , n73975 );
or ( n73977 , n73973 , n73897 );
nand ( n73978 , n73976 , n73977 );
and ( n73979 , n73978 , n73909 );
and ( n73980 , n72452 , n69359 );
nor ( n73981 , n73979 , n73980 );
or ( n73982 , n73981 , n70210 );
nor ( n73983 , n72633 , n72626 );
not ( n73984 , n73983 );
not ( n73985 , n73916 );
not ( n73986 , n69743 );
or ( n73987 , n73985 , n73986 );
or ( n73988 , n69743 , n73916 );
nand ( n73989 , n73987 , n73988 );
not ( n73990 , n73989 );
or ( n73991 , n73984 , n73990 );
or ( n73992 , n73983 , n73989 );
nand ( n73993 , n73991 , n73992 );
not ( n73994 , n73993 );
nor ( n73995 , n72570 , n72638 );
not ( n73996 , n73995 );
nor ( n73997 , n73996 , n72522 );
not ( n73998 , n73997 );
not ( n73999 , n70553 );
or ( n74000 , n73998 , n73999 );
not ( n74001 , n73995 );
not ( n74002 , n72604 );
or ( n74003 , n74001 , n74002 );
not ( n74004 , n72639 );
not ( n74005 , n72620 );
or ( n74006 , n74004 , n74005 );
nand ( n74007 , n74006 , n72640 );
not ( n74008 , n74007 );
nand ( n74009 , n74003 , n74008 );
not ( n74010 , n74009 );
nand ( n74011 , n74000 , n74010 );
not ( n74012 , n74011 );
or ( n74013 , n73994 , n74012 );
or ( n74014 , n74011 , n73993 );
nand ( n74015 , n74013 , n74014 );
nand ( n74016 , n74015 , n70568 );
xor ( n74017 , n73916 , n69743 );
not ( n74018 , n74017 );
and ( n74019 , n72626 , n69729 );
not ( n74020 , n74019 );
or ( n74021 , n74018 , n74020 );
or ( n74022 , n74019 , n74017 );
nand ( n74023 , n74021 , n74022 );
not ( n74024 , n74023 );
nand ( n74025 , n72674 , n72771 );
nor ( n74026 , n74025 , n72724 );
not ( n74027 , n74026 );
not ( n74028 , n70809 );
or ( n74029 , n74027 , n74028 );
not ( n74030 , n72749 );
not ( n74031 , n74025 );
and ( n74032 , n74030 , n74031 );
not ( n74033 , n72771 );
not ( n74034 , n72766 );
or ( n74035 , n74033 , n74034 );
nand ( n74036 , n74035 , n72772 );
nor ( n74037 , n74032 , n74036 );
nand ( n74038 , n74029 , n74037 );
not ( n74039 , n74038 );
or ( n74040 , n74024 , n74039 );
or ( n74041 , n74038 , n74023 );
nand ( n74042 , n74040 , n74041 );
and ( n74043 , n74042 , n70573 );
nand ( n74044 , n72797 , n70876 , n69721 );
not ( n74045 , n73916 );
not ( n74046 , n72626 );
nand ( n74047 , n74046 , n72812 , n72817 );
nor ( n74048 , n70832 , n74047 );
not ( n74049 , n74048 );
or ( n74050 , n74045 , n74049 );
or ( n74051 , n74048 , n73916 );
nand ( n74052 , n74050 , n74051 );
nand ( n74053 , n74052 , n73766 );
nand ( n74054 , n70849 , n73916 );
nand ( n74055 , n70870 , n69741 );
nand ( n74056 , n74044 , n74053 , n74054 , n74055 );
nor ( n74057 , n74043 , n74056 );
nand ( n74058 , n73982 , n74016 , n74057 );
buf ( n7920 , n74058 );
buf ( n7921 , 1'b0 );
not ( n74061 , n68838 );
buf ( n74062 , n74061 );
buf ( n74063 , n68634 );
or ( n74064 , n72470 , n70210 );
nand ( n74065 , n72646 , n70568 );
and ( n74066 , n72778 , n70573 );
nand ( n74067 , n72801 , n70876 );
nand ( n74068 , n72823 , n70840 );
nand ( n74069 , n70849 , n72626 );
nand ( n74070 , n70870 , n69710 );
nand ( n74071 , n74067 , n74068 , n74069 , n74070 );
nor ( n74072 , n74066 , n74071 );
and ( n74073 , n74065 , n74072 );
nand ( n74074 , n74064 , n74073 );
buf ( n7936 , n74074 );
buf ( n7937 , 1'b0 );
not ( n74077 , n68838 );
buf ( n74078 , n74077 );
buf ( n74079 , n68634 );
or ( n74080 , n72845 , n70210 );
nand ( n74081 , n72866 , n70568 );
and ( n74082 , n72889 , n70573 );
not ( n74083 , n72894 );
nand ( n74084 , n74083 , n70876 );
nand ( n74085 , n72906 , n73766 );
nand ( n74086 , n70849 , n72815 );
nand ( n74087 , n70870 , n69688 );
nand ( n74088 , n74084 , n74085 , n74086 , n74087 );
nor ( n74089 , n74082 , n74088 );
and ( n74090 , n74081 , n74089 );
nand ( n74091 , n74080 , n74090 );
buf ( n7953 , n74091 );
buf ( n74093 , 1'b0 );
not ( n74094 , n68838 );
buf ( n74095 , n74094 );
buf ( n74096 , n68634 );
or ( n74097 , n72933 , n70210 );
nand ( n74098 , n72952 , n70568 );
and ( n74099 , n72967 , n70573 );
nor ( n74100 , n72972 , n73863 );
not ( n74101 , n72534 );
nor ( n74102 , n74101 , n70848 );
nor ( n74103 , n74100 , n74102 );
nand ( n74104 , n72982 , n70840 );
nand ( n74105 , n70870 , n69670 );
nand ( n74106 , n74103 , n74104 , n74105 );
nor ( n74107 , n74099 , n74106 );
and ( n74108 , n74098 , n74107 );
nand ( n74109 , n74097 , n74108 );
buf ( n7971 , n74109 );
buf ( n7972 , 1'b0 );
not ( n74112 , n68838 );
buf ( n74113 , n74112 );
buf ( n74114 , n68634 );
or ( n74115 , n73007 , n70210 );
nand ( n74116 , n73022 , n70568 );
and ( n74117 , n73040 , n70573 );
nand ( n74118 , n73056 , n73766 );
and ( n74119 , n70849 , n72544 );
nor ( n74120 , n73045 , n73863 );
nor ( n74121 , n74119 , n74120 );
nand ( n74122 , n70870 , n69831 );
nand ( n74123 , n74118 , n74121 , n74122 );
nor ( n74124 , n74117 , n74123 );
and ( n74125 , n74116 , n74124 );
nand ( n74126 , n74115 , n74125 );
buf ( n7988 , n74126 );
buf ( n7989 , 1'b0 );
not ( n74129 , n68838 );
buf ( n74130 , n74129 );
buf ( n7992 , n68634 );
or ( n74132 , n73079 , n70210 );
nand ( n74133 , n73092 , n70568 );
and ( n74134 , n73104 , n70573 );
nand ( n74135 , n73117 , n73766 );
not ( n74136 , n73109 );
not ( n74137 , n70875 );
and ( n74138 , n74136 , n74137 );
and ( n74139 , n70849 , n72557 );
nor ( n74140 , n74138 , n74139 );
nand ( n74141 , n70870 , n69916 );
nand ( n74142 , n74135 , n74140 , n74141 );
nor ( n74143 , n74134 , n74142 );
and ( n74144 , n74133 , n74143 );
nand ( n74145 , n74132 , n74144 );
buf ( n74146 , n74145 );
buf ( n74147 , 1'b0 );
not ( n74148 , n68838 );
buf ( n8010 , n74148 );
buf ( n8011 , n68634 );
or ( n74151 , n73143 , n70210 );
nand ( n74152 , n73161 , n70568 );
and ( n74153 , n73189 , n70573 );
nand ( n74154 , n73202 , n73766 );
not ( n74155 , n73194 );
not ( n74156 , n70875 );
and ( n74157 , n74155 , n74156 );
and ( n74158 , n70849 , n72510 );
nor ( n74159 , n74157 , n74158 );
nand ( n74160 , n70870 , n69749 );
nand ( n74161 , n74154 , n74159 , n74160 );
nor ( n74162 , n74153 , n74161 );
and ( n74163 , n74152 , n74162 );
nand ( n74164 , n74151 , n74163 );
buf ( n8026 , n74164 );
buf ( n8027 , 1'b0 );
not ( n74167 , n68838 );
buf ( n74168 , n74167 );
buf ( n74169 , n68634 );
or ( n74170 , n73224 , n70210 );
nand ( n74171 , n73239 , n70568 );
and ( n74172 , n73253 , n70573 );
nand ( n74173 , n73266 , n73766 );
not ( n74174 , n73258 );
not ( n74175 , n70875 );
and ( n74176 , n74174 , n74175 );
and ( n74177 , n70849 , n72499 );
nor ( n74178 , n74176 , n74177 );
nand ( n74179 , n70870 , n69783 );
nand ( n74180 , n74173 , n74178 , n74179 );
nor ( n74181 , n74172 , n74180 );
and ( n74182 , n74171 , n74181 );
nand ( n74183 , n74170 , n74182 );
buf ( n8045 , n74183 );
buf ( n8046 , 1'b0 );
not ( n74186 , n68838 );
buf ( n74187 , n74186 );
buf ( n74188 , n68634 );
or ( n74189 , n73289 , n70210 );
nand ( n74190 , n73304 , n70568 );
and ( n74191 , n73323 , n70573 );
nand ( n74192 , n73337 , n73766 );
not ( n74193 , n70875 );
not ( n74194 , n73328 );
and ( n74195 , n74193 , n74194 );
and ( n74196 , n70849 , n72475 );
nor ( n74197 , n74195 , n74196 );
nand ( n74198 , n70870 , n69876 );
nand ( n74199 , n74192 , n74197 , n74198 );
nor ( n74200 , n74191 , n74199 );
and ( n74201 , n74190 , n74200 );
nand ( n74202 , n74189 , n74201 );
buf ( n74203 , n74202 );
buf ( n74204 , 1'b0 );
not ( n74205 , n68838 );
buf ( n8067 , n74205 );
buf ( n8068 , n68634 );
or ( n74208 , n73361 , n70210 );
nand ( n74209 , n73369 , n70568 );
and ( n74210 , n70573 , n73381 );
nand ( n74211 , n73394 , n73766 );
not ( n74212 , n70875 );
not ( n74213 , n73386 );
and ( n74214 , n74212 , n74213 );
and ( n74215 , n70849 , n72485 );
nor ( n74216 , n74214 , n74215 );
nand ( n74217 , n70870 , n69862 );
nand ( n74218 , n74211 , n74216 , n74217 );
nor ( n74219 , n74210 , n74218 );
and ( n74220 , n74209 , n74219 );
nand ( n74221 , n74208 , n74220 );
buf ( n74222 , n74221 );
buf ( n8084 , 1'b0 );
not ( n74224 , n68838 );
buf ( n74225 , n74224 );
buf ( n74226 , n68634 );
or ( n74227 , n73416 , n70210 );
not ( n74228 , n73435 );
or ( n74229 , n73765 , n74228 );
not ( n74230 , n70051 );
or ( n74231 , n73843 , n74230 );
not ( n74232 , n70503 );
or ( n74233 , n70848 , n74232 );
nand ( n74234 , n74229 , n74231 , n74233 );
not ( n74235 , n73426 );
not ( n74236 , n70568 );
or ( n74237 , n74235 , n74236 );
nand ( n74238 , n70573 , n73428 );
nand ( n74239 , n70876 , n70041 );
nand ( n74240 , n74237 , n74238 , n74239 );
nor ( n74241 , n74234 , n74240 );
nand ( n74242 , n74227 , n74241 );
buf ( n74243 , n74242 );
buf ( n74244 , 1'b0 );
not ( n74245 , n68838 );
buf ( n74246 , n74245 );
buf ( n74247 , n68634 );
or ( n74248 , n73445 , n70210 );
nand ( n74249 , n71134 , n70568 );
and ( n74250 , n71188 , n70573 );
nand ( n74251 , n71200 , n73766 );
not ( n74252 , n70875 );
not ( n74253 , n73453 );
and ( n74254 , n74252 , n74253 );
and ( n74255 , n70849 , n71122 );
nor ( n74256 , n74254 , n74255 );
nand ( n74257 , n70870 , n69798 );
nand ( n74258 , n74251 , n74256 , n74257 );
nor ( n74259 , n74250 , n74258 );
and ( n74260 , n74249 , n74259 );
nand ( n74261 , n74248 , n74260 );
buf ( n74262 , n74261 );
buf ( n74263 , 1'b0 );
not ( n74264 , n68838 );
buf ( n8126 , n74264 );
buf ( n8127 , n68634 );
or ( n74267 , n73468 , n70210 );
nand ( n74268 , n71233 , n70568 );
and ( n74269 , n71248 , n70573 );
nand ( n74270 , n71256 , n70840 );
not ( n74271 , n70875 );
not ( n74272 , n73475 );
and ( n74273 , n74271 , n74272 );
and ( n74274 , n70849 , n71092 );
nor ( n74275 , n74273 , n74274 );
nand ( n74276 , n70870 , n69806 );
nand ( n74277 , n74270 , n74275 , n74276 );
nor ( n74278 , n74269 , n74277 );
and ( n74279 , n74268 , n74278 );
nand ( n74280 , n74267 , n74279 );
buf ( n8142 , n74280 );
buf ( n8143 , 1'b0 );
not ( n74283 , n68838 );
buf ( n74284 , n74283 );
buf ( n74285 , n68634 );
or ( n74286 , n71281 , n70210 );
nand ( n74287 , n71291 , n70568 );
and ( n74288 , n71304 , n70573 );
nand ( n74289 , n71312 , n70840 );
not ( n74290 , n70875 );
not ( n74291 , n73497 );
and ( n74292 , n74290 , n74291 );
and ( n74293 , n70849 , n71074 );
nor ( n74294 , n74292 , n74293 );
nand ( n74295 , n73844 , n69651 );
nand ( n74296 , n74289 , n74294 , n74295 );
nor ( n74297 , n74288 , n74296 );
nand ( n74298 , n74286 , n74287 , n74297 );
buf ( n74299 , n74298 );
buf ( n74300 , 1'b0 );
not ( n74301 , n68838 );
buf ( n8163 , n74301 );
buf ( n8164 , n68634 );
or ( n74304 , n73532 , n70210 );
and ( n74305 , n70573 , n71416 );
nand ( n74306 , n71428 , n70840 );
not ( n74307 , n73863 );
not ( n74308 , n73539 );
and ( n74309 , n74307 , n74308 );
and ( n74310 , n70849 , n70238 );
nor ( n74311 , n74309 , n74310 );
nand ( n74312 , n73844 , n3466 );
nand ( n74313 , n74306 , n74311 , n74312 );
nor ( n74314 , n74305 , n74313 );
nand ( n74315 , n71390 , n70568 );
and ( n74316 , n74314 , n74315 );
nand ( n74317 , n74304 , n74316 );
buf ( n74318 , n74317 );
buf ( n74319 , 1'b0 );
not ( n74320 , n68838 );
buf ( n74321 , n74320 );
buf ( n74322 , n68634 );
or ( n74323 , n73557 , n70210 );
and ( n74324 , n70573 , n71491 );
nand ( n74325 , n71501 , n73766 );
not ( n74326 , n70875 );
not ( n74327 , n73563 );
and ( n74328 , n74326 , n74327 );
and ( n74329 , n70849 , n70327 );
nor ( n74330 , n74328 , n74329 );
nand ( n74331 , n73844 , n3450 );
nand ( n74332 , n74325 , n74330 , n74331 );
nor ( n74333 , n74324 , n74332 );
nand ( n74334 , n71475 , n70568 );
and ( n74335 , n74333 , n74334 );
nand ( n74336 , n74323 , n74335 );
buf ( n74337 , n74336 );
buf ( n8199 , 1'b0 );
not ( n74339 , n68838 );
buf ( n8201 , n74339 );
buf ( n8202 , n68634 );
or ( n74342 , n73591 , n70210 );
and ( n74343 , n70573 , n73633 );
nand ( n74344 , n73642 , n70840 );
not ( n74345 , n70875 );
not ( n74346 , n73598 );
and ( n74347 , n74345 , n74346 );
and ( n74348 , n70849 , n70296 );
nor ( n74349 , n74347 , n74348 );
nand ( n74350 , n73844 , n69558 );
nand ( n74351 , n74344 , n74349 , n74350 );
nor ( n74352 , n74343 , n74351 );
nand ( n74353 , n73614 , n70568 );
and ( n74354 , n74352 , n74353 );
nand ( n74355 , n74342 , n74354 );
buf ( n8217 , n74355 );
buf ( n74357 , 1'b0 );
not ( n74358 , n68838 );
buf ( n74359 , n74358 );
buf ( n8221 , n68634 );
or ( n74361 , n73655 , n70210 );
and ( n74362 , n70573 , n71558 );
nand ( n74363 , n71567 , n73766 );
not ( n74364 , n70875 );
not ( n74365 , n73662 );
and ( n74366 , n74364 , n74365 );
and ( n74367 , n70849 , n70308 );
nor ( n74368 , n74366 , n74367 );
nand ( n74369 , n73844 , n69577 );
nand ( n74370 , n74363 , n74368 , n74369 );
nor ( n74371 , n74362 , n74370 );
nand ( n74372 , n71545 , n70568 );
and ( n74373 , n74371 , n74372 );
nand ( n74374 , n74361 , n74373 );
buf ( n74375 , n74374 );
buf ( n8237 , 1'b0 );
not ( n74377 , n68838 );
buf ( n74378 , n74377 );
buf ( n74379 , n68634 );
or ( n74380 , n73680 , n70210 );
and ( n74381 , n70573 , n71638 );
nand ( n74382 , n71647 , n70840 );
not ( n74383 , n70875 );
not ( n74384 , n73686 );
and ( n74385 , n74383 , n74384 );
and ( n74386 , n70849 , n70273 );
nor ( n74387 , n74385 , n74386 );
nand ( n74388 , n73844 , n69507 );
nand ( n74389 , n74382 , n74387 , n74388 );
nor ( n74390 , n74381 , n74389 );
nand ( n74391 , n71618 , n70568 );
and ( n74392 , n74390 , n74391 );
nand ( n74393 , n74380 , n74392 );
buf ( n74394 , n74393 );
buf ( n74395 , 1'b0 );
not ( n74396 , n68838 );
buf ( n74397 , n74396 );
buf ( n74398 , n68634 );
or ( n74399 , n73704 , n70210 );
and ( n74400 , n70573 , n71699 );
nand ( n74401 , n71707 , n70840 );
not ( n74402 , n73863 );
not ( n74403 , n73711 );
and ( n74404 , n74402 , n74403 );
and ( n74405 , n70849 , n70253 );
nor ( n74406 , n74404 , n74405 );
nand ( n74407 , n73844 , n69522 );
nand ( n74408 , n74401 , n74406 , n74407 );
nor ( n74409 , n74400 , n74408 );
nand ( n74410 , n71685 , n70568 );
and ( n74411 , n74409 , n74410 );
nand ( n74412 , n74399 , n74411 );
buf ( n8274 , n74412 );
buf ( n8275 , 1'b0 );
not ( n74415 , n68838 );
buf ( n8277 , n74415 );
buf ( n74417 , n68634 );
or ( n74418 , n73735 , n70210 );
not ( n74419 , n3815 );
not ( n74420 , n70870 );
or ( n74421 , n74419 , n74420 );
or ( n74422 , n70840 , n70849 );
nand ( n74423 , n74422 , n70522 );
nand ( n74424 , n74421 , n74423 );
nand ( n74425 , n70568 , n73745 );
nand ( n74426 , n70573 , n73753 );
nand ( n74427 , n70876 , n69950 );
nand ( n74428 , n74425 , n74426 , n74427 );
nor ( n74429 , n74424 , n74428 );
nand ( n74430 , n74418 , n74429 );
buf ( n74431 , n74430 );
buf ( n74432 , 1'b0 );
not ( n74433 , n68838 );
buf ( n8295 , n74433 );
buf ( n8296 , n68634 );
and ( n74436 , n72040 , n70196 );
nand ( n74437 , n72055 , n70929 );
nand ( n74438 , n72048 , n70571 );
not ( n74439 , n73794 );
not ( n74440 , n70846 );
and ( n74441 , n74439 , n74440 );
and ( n74442 , n72069 , n70995 );
nor ( n74443 , n74441 , n74442 );
nand ( n74444 , n74437 , n74438 , n74443 );
nor ( n74445 , n74436 , n74444 );
or ( n74446 , n74445 , n71016 );
nand ( n74447 , n71016 , n69546 );
nand ( n74448 , n74446 , n74447 );
buf ( n74449 , n74448 );
buf ( n8311 , 1'b0 );
not ( n74451 , n68838 );
buf ( n74452 , n74451 );
buf ( n74453 , n68634 );
not ( n74454 , n72094 );
and ( n74455 , n74454 , n70923 );
not ( n74456 , n70929 );
not ( n74457 , n72112 );
or ( n74458 , n74456 , n74457 );
and ( n74459 , n72130 , n70571 );
not ( n74460 , n70847 );
not ( n74461 , n70388 );
or ( n74462 , n74460 , n74461 );
nand ( n74463 , n72150 , n70995 );
nand ( n74464 , n74462 , n74463 );
nor ( n74465 , n74459 , n74464 );
nand ( n74466 , n74458 , n74465 );
nor ( n74467 , n74455 , n74466 );
or ( n74468 , n74467 , n71016 );
not ( n74469 , n71016 );
not ( n74470 , n74469 );
nand ( n74471 , n74470 , n3316 );
nand ( n74472 , n74468 , n74471 );
buf ( n74473 , n74472 );
buf ( n74474 , 1'b0 );
not ( n74475 , n68838 );
buf ( n74476 , n74475 );
buf ( n74477 , n68634 );
not ( n74478 , n72169 );
and ( n74479 , n74478 , n70923 );
nand ( n74480 , n72191 , n70931 );
nand ( n74481 , n72178 , n70571 );
and ( n74482 , n70477 , n70847 );
and ( n74483 , n72207 , n70995 );
nor ( n74484 , n74482 , n74483 );
nand ( n74485 , n74480 , n74481 , n74484 );
nor ( n74486 , n74479 , n74485 );
or ( n74487 , n74486 , n71016 );
not ( n74488 , n71343 );
nand ( n74489 , n74488 , n3282 );
nand ( n74490 , n74487 , n74489 );
buf ( n74491 , n74490 );
buf ( n8353 , 1'b0 );
not ( n74493 , n68838 );
buf ( n74494 , n74493 );
buf ( n74495 , n68634 );
not ( n74496 , n72230 );
and ( n74497 , n74496 , n70923 );
not ( n74498 , n70929 );
not ( n74499 , n72242 );
or ( n74500 , n74498 , n74499 );
and ( n74501 , n72254 , n70571 );
not ( n74502 , n70847 );
not ( n74503 , n70432 );
or ( n74504 , n74502 , n74503 );
nand ( n74505 , n72269 , n70995 );
nand ( n74506 , n74504 , n74505 );
nor ( n74507 , n74501 , n74506 );
nand ( n74508 , n74500 , n74507 );
nor ( n74509 , n74497 , n74508 );
or ( n74510 , n74509 , n71016 );
nand ( n74511 , n74470 , n69492 );
nand ( n74512 , n74510 , n74511 );
buf ( n74513 , n74512 );
buf ( n74514 , 1'b0 );
not ( n74515 , n68838 );
buf ( n74516 , n74515 );
buf ( n74517 , n68634 );
and ( n74518 , n72289 , n70923 );
not ( n74519 , n70929 );
not ( n74520 , n72293 );
or ( n74521 , n74519 , n74520 );
and ( n74522 , n72300 , n70571 );
not ( n74523 , n72302 );
not ( n74524 , n70847 );
or ( n74525 , n74523 , n74524 );
not ( n74526 , n70995 );
or ( n74527 , n73867 , n74526 );
nand ( n74528 , n74525 , n74527 );
nor ( n74529 , n74522 , n74528 );
nand ( n74530 , n74521 , n74529 );
nor ( n74531 , n74518 , n74530 );
or ( n74532 , n74531 , n71344 );
nand ( n74533 , n74488 , n3342 );
nand ( n74534 , n74532 , n74533 );
buf ( n8396 , n74534 );
buf ( n8397 , 1'b0 );
not ( n74537 , n68838 );
buf ( n74538 , n74537 );
buf ( n74539 , n68634 );
not ( n74540 , n74469 );
or ( n74541 , n72340 , n70195 );
and ( n74542 , n72356 , n70571 );
not ( n74543 , n70420 );
not ( n74544 , n70847 );
or ( n74545 , n74543 , n74544 );
nand ( n74546 , n72365 , n70995 );
nand ( n74547 , n74545 , n74546 );
nor ( n74548 , n74542 , n74547 );
nand ( n74549 , n72345 , n70929 );
and ( n74550 , n74548 , n74549 );
nand ( n74551 , n74541 , n74550 );
not ( n74552 , n74551 );
or ( n74553 , n74540 , n74552 );
nand ( n74554 , n71344 , n3301 );
nand ( n74555 , n74553 , n74554 );
buf ( n8417 , n74555 );
buf ( n74557 , 1'b0 );
not ( n74558 , n68838 );
buf ( n74559 , n74558 );
buf ( n8421 , n68634 );
and ( n74561 , n71016 , n69936 );
not ( n74562 , n71016 );
and ( n74563 , n74562 , n73928 );
or ( n74564 , n74561 , n74563 );
buf ( n74565 , n74564 );
buf ( n8427 , 1'b0 );
not ( n74567 , n68838 );
buf ( n74568 , n74567 );
buf ( n74569 , n68634 );
not ( n74570 , n73948 );
or ( n74571 , n74570 , n74470 );
or ( n74572 , n71343 , n69898 );
nand ( n74573 , n74571 , n74572 );
buf ( n74574 , n74573 );
buf ( n8436 , 1'b0 );
not ( n74576 , n68838 );
buf ( n8438 , n74576 );
buf ( n8439 , n68634 );
not ( n74579 , n72384 );
and ( n74580 , n74579 , n70196 );
not ( n74581 , n70929 );
not ( n74582 , n72405 );
or ( n74583 , n74581 , n74582 );
and ( n74584 , n72418 , n70571 );
or ( n74585 , n72410 , n70846 );
or ( n74586 , n72394 , n74526 );
nand ( n74587 , n74585 , n74586 );
nor ( n74588 , n74584 , n74587 );
nand ( n74589 , n74583 , n74588 );
nor ( n74590 , n74580 , n74589 );
or ( n74591 , n74590 , n71016 );
nand ( n74592 , n71344 , n70069 );
nand ( n74593 , n74591 , n74592 );
buf ( n8455 , n74593 );
buf ( n74595 , 1'b0 );
not ( n74596 , n68838 );
buf ( n74597 , n74596 );
buf ( n8459 , n68634 );
not ( n74599 , n73981 );
and ( n74600 , n74599 , n70196 );
not ( n74601 , n70929 );
not ( n74602 , n74015 );
or ( n74603 , n74601 , n74602 );
and ( n74604 , n74042 , n70571 );
not ( n74605 , n70995 );
not ( n74606 , n74052 );
or ( n74607 , n74605 , n74606 );
nand ( n74608 , n70847 , n73916 );
nand ( n74609 , n74607 , n74608 );
nor ( n74610 , n74604 , n74609 );
nand ( n74611 , n74603 , n74610 );
nor ( n74612 , n74600 , n74611 );
or ( n74613 , n74612 , n74488 );
nand ( n74614 , n71344 , n69737 );
nand ( n74615 , n74613 , n74614 );
buf ( n74616 , n74615 );
buf ( n74617 , 1'b0 );
not ( n74618 , n68838 );
buf ( n74619 , n74618 );
buf ( n74620 , n68634 );
not ( n74621 , n72470 );
not ( n74622 , n70923 );
not ( n74623 , n74622 );
and ( n74624 , n74621 , n74623 );
nand ( n74625 , n72646 , n70929 );
and ( n74626 , n72778 , n70571 );
not ( n74627 , n70995 );
not ( n74628 , n72823 );
or ( n74629 , n74627 , n74628 );
nand ( n74630 , n70847 , n72626 );
nand ( n74631 , n74629 , n74630 );
nor ( n74632 , n74626 , n74631 );
nand ( n74633 , n74625 , n74632 );
nor ( n74634 , n74624 , n74633 );
or ( n74635 , n74634 , n74488 );
nand ( n74636 , n74470 , n69715 );
nand ( n74637 , n74635 , n74636 );
buf ( n8499 , n74637 );
buf ( n74639 , 1'b0 );
not ( n74640 , n68838 );
buf ( n8502 , n74640 );
buf ( n74642 , n68634 );
not ( n74643 , n72845 );
and ( n74644 , n74643 , n74623 );
and ( n74645 , n72889 , n70571 );
not ( n74646 , n70995 );
not ( n74647 , n72906 );
or ( n74648 , n74646 , n74647 );
nand ( n74649 , n70847 , n72815 );
nand ( n74650 , n74648 , n74649 );
nor ( n74651 , n74645 , n74650 );
nand ( n74652 , n72866 , n70929 );
nand ( n74653 , n74651 , n74652 );
nor ( n74654 , n74644 , n74653 );
or ( n74655 , n74654 , n74488 );
nand ( n74656 , n74470 , n69693 );
nand ( n74657 , n74655 , n74656 );
buf ( n8519 , n74657 );
buf ( n8520 , 1'b0 );
not ( n74660 , n68838 );
buf ( n74661 , n74660 );
buf ( n74662 , n68634 );
not ( n74663 , n72933 );
and ( n74664 , n74663 , n70196 );
nand ( n74665 , n72952 , n70929 );
and ( n74666 , n72967 , n70571 );
not ( n74667 , n70995 );
not ( n74668 , n72982 );
or ( n74669 , n74667 , n74668 );
nand ( n74670 , n70847 , n72534 );
nand ( n74671 , n74669 , n74670 );
nor ( n74672 , n74666 , n74671 );
nand ( n74673 , n74665 , n74672 );
nor ( n74674 , n74664 , n74673 );
or ( n74675 , n74674 , n71016 );
nand ( n74676 , n71344 , n69665 );
nand ( n74677 , n74675 , n74676 );
buf ( n8539 , n74677 );
buf ( n8540 , 1'b0 );
not ( n74680 , n68838 );
buf ( n74681 , n74680 );
buf ( n74682 , n68634 );
not ( n74683 , n73007 );
and ( n74684 , n74683 , n74623 );
nand ( n74685 , n73022 , n70929 );
and ( n74686 , n70571 , n73040 );
not ( n74687 , n70995 );
not ( n74688 , n73056 );
or ( n74689 , n74687 , n74688 );
nand ( n74690 , n70847 , n72544 );
nand ( n74691 , n74689 , n74690 );
nor ( n74692 , n74686 , n74691 );
nand ( n74693 , n74685 , n74692 );
nor ( n74694 , n74684 , n74693 );
or ( n74695 , n74694 , n71344 );
nand ( n74696 , n74470 , n69837 );
nand ( n74697 , n74695 , n74696 );
buf ( n74698 , n74697 );
buf ( n74699 , 1'b0 );
not ( n74700 , n68838 );
buf ( n74701 , n74700 );
buf ( n8563 , n68634 );
not ( n74703 , n73079 );
and ( n74704 , n74703 , n70923 );
nand ( n74705 , n73092 , n70929 );
and ( n74706 , n73104 , n70571 );
not ( n74707 , n70995 );
not ( n74708 , n73117 );
or ( n74709 , n74707 , n74708 );
nand ( n74710 , n70847 , n72557 );
nand ( n74711 , n74709 , n74710 );
nor ( n74712 , n74706 , n74711 );
nand ( n74713 , n74705 , n74712 );
nor ( n74714 , n74704 , n74713 );
or ( n74715 , n74714 , n74470 );
nand ( n74716 , n74470 , n69912 );
nand ( n74717 , n74715 , n74716 );
buf ( n74718 , n74717 );
buf ( n8580 , 1'b0 );
not ( n74720 , n68838 );
buf ( n74721 , n74720 );
buf ( n74722 , n68634 );
not ( n74723 , n73143 );
and ( n74724 , n74723 , n70923 );
nand ( n74725 , n73161 , n70929 );
and ( n74726 , n73189 , n70571 );
not ( n74727 , n70995 );
not ( n74728 , n73202 );
or ( n74729 , n74727 , n74728 );
nand ( n74730 , n70847 , n72510 );
nand ( n74731 , n74729 , n74730 );
nor ( n74732 , n74726 , n74731 );
nand ( n74733 , n74725 , n74732 );
nor ( n74734 , n74724 , n74733 );
or ( n74735 , n74734 , n71344 );
nand ( n74736 , n74488 , n69755 );
nand ( n74737 , n74735 , n74736 );
buf ( n74738 , n74737 );
buf ( n74739 , 1'b0 );
not ( n74740 , n68838 );
buf ( n8602 , n74740 );
buf ( n8603 , n68634 );
not ( n74743 , n73224 );
and ( n74744 , n74743 , n70923 );
nand ( n74745 , n73239 , n70929 );
and ( n74746 , n73253 , n70571 );
not ( n74747 , n70995 );
not ( n74748 , n73266 );
or ( n74749 , n74747 , n74748 );
nand ( n74750 , n70847 , n72499 );
nand ( n74751 , n74749 , n74750 );
nor ( n74752 , n74746 , n74751 );
nand ( n74753 , n74745 , n74752 );
nor ( n74754 , n74744 , n74753 );
or ( n74755 , n74754 , n71344 );
nand ( n74756 , n74488 , n69777 );
nand ( n74757 , n74755 , n74756 );
buf ( n8619 , n74757 );
buf ( n74759 , 1'b0 );
not ( n74760 , n68838 );
buf ( n74761 , n74760 );
buf ( n74762 , n68634 );
not ( n74763 , n73289 );
and ( n74764 , n74763 , n70923 );
nand ( n74765 , n73304 , n70929 );
and ( n74766 , n73323 , n70571 );
not ( n74767 , n70995 );
not ( n74768 , n73337 );
or ( n74769 , n74767 , n74768 );
nand ( n74770 , n70847 , n72475 );
nand ( n74771 , n74769 , n74770 );
nor ( n74772 , n74766 , n74771 );
nand ( n74773 , n74765 , n74772 );
nor ( n74774 , n74764 , n74773 );
or ( n74775 , n74774 , n74470 );
nand ( n74776 , n74488 , n69882 );
nand ( n74777 , n74775 , n74776 );
buf ( n8639 , n74777 );
buf ( n74779 , 1'b0 );
not ( n74780 , n68838 );
buf ( n74781 , n74780 );
buf ( n8643 , n68634 );
not ( n74783 , n73361 );
and ( n74784 , n74783 , n74623 );
not ( n74785 , n70929 );
not ( n74786 , n73369 );
or ( n74787 , n74785 , n74786 );
and ( n74788 , n73381 , n70571 );
not ( n74789 , n70995 );
not ( n74790 , n73394 );
or ( n74791 , n74789 , n74790 );
nand ( n74792 , n70847 , n72485 );
nand ( n74793 , n74791 , n74792 );
nor ( n74794 , n74788 , n74793 );
nand ( n74795 , n74787 , n74794 );
nor ( n74796 , n74784 , n74795 );
or ( n74797 , n74796 , n71344 );
nand ( n74798 , n74470 , n69856 );
nand ( n74799 , n74797 , n74798 );
buf ( n8661 , n74799 );
buf ( n74801 , 1'b0 );
not ( n74802 , n68838 );
buf ( n74803 , n74802 );
buf ( n8665 , n68634 );
not ( n74805 , n73416 );
and ( n74806 , n74805 , n70196 );
not ( n74807 , n70929 );
not ( n74808 , n73426 );
or ( n74809 , n74807 , n74808 );
and ( n74810 , n73428 , n70571 );
and ( n74811 , n70847 , n70503 );
and ( n74812 , n73435 , n70995 );
nor ( n74813 , n74810 , n74811 , n74812 );
nand ( n74814 , n74809 , n74813 );
nor ( n74815 , n74806 , n74814 );
or ( n74816 , n74815 , n71016 );
nand ( n74817 , n71344 , n70049 );
nand ( n74818 , n74816 , n74817 );
buf ( n74819 , n74818 );
buf ( n8681 , 1'b0 );
not ( n74821 , n68838 );
buf ( n74822 , n74821 );
buf ( n74823 , n68634 );
and ( n74824 , n73590 , n70923 );
not ( n74825 , n70931 );
not ( n74826 , n73614 );
or ( n74827 , n74825 , n74826 );
and ( n74828 , n73633 , n70571 );
not ( n74829 , n70995 );
not ( n74830 , n73642 );
or ( n74831 , n74829 , n74830 );
nand ( n74832 , n70296 , n70847 );
nand ( n74833 , n74831 , n74832 );
nor ( n74834 , n74828 , n74833 );
nand ( n74835 , n74827 , n74834 );
nor ( n74836 , n74824 , n74835 );
or ( n74837 , n74836 , n71016 );
nand ( n74838 , n71016 , n69562 );
nand ( n74839 , n74837 , n74838 );
buf ( n74840 , n74839 );
buf ( n74841 , 1'b0 );
not ( n74842 , n68838 );
buf ( n74843 , n74842 );
buf ( n74844 , n68634 );
not ( n74845 , n73735 );
not ( n74846 , n70195 );
and ( n74847 , n74845 , n74846 );
not ( n74848 , n70571 );
not ( n74849 , n73753 );
or ( n74850 , n74848 , n74849 );
and ( n74851 , n73745 , n70929 );
nand ( n74852 , n70846 , n74526 );
and ( n74853 , n74852 , n70522 );
nor ( n74854 , n74851 , n74853 );
nand ( n74855 , n74850 , n74854 );
nor ( n74856 , n74847 , n74855 );
or ( n74857 , n74856 , n71016 );
nand ( n74858 , n71016 , n69957 );
nand ( n74859 , n74857 , n74858 );
buf ( n8721 , n74859 );
buf ( n74861 , 1'b0 );
not ( n74862 , n68838 );
buf ( n8724 , n74862 );
buf ( n74864 , n68634 );
not ( n74865 , n70164 );
and ( n74866 , n70148 , n74865 , n70181 , n70854 );
not ( n74867 , n74866 );
or ( n74868 , n71015 , n74867 );
nand ( n74869 , n74867 , n69541 );
nand ( n74870 , n74868 , n74869 );
buf ( n8732 , n74870 );
buf ( n8733 , 1'b0 );
not ( n74873 , n68838 );
buf ( n8735 , n74873 );
buf ( n74875 , n68634 );
or ( n74876 , n74445 , n74867 );
nand ( n74877 , n74867 , n3412 );
nand ( n74878 , n74876 , n74877 );
buf ( n8740 , n74878 );
buf ( n8741 , 1'b0 );
not ( n74881 , n68838 );
buf ( n74882 , n74881 );
buf ( n74883 , n68634 );
or ( n74884 , n74467 , n74867 );
nand ( n74885 , n74867 , n69468 );
nand ( n74886 , n74884 , n74885 );
buf ( n74887 , n74886 );
buf ( n74888 , 1'b0 );
not ( n74889 , n68838 );
buf ( n8751 , n74889 );
buf ( n74891 , n68634 );
or ( n74892 , n74486 , n74867 );
nand ( n74893 , n74867 , n69433 );
nand ( n74894 , n74892 , n74893 );
buf ( n8756 , n74894 );
buf ( n74896 , 1'b0 );
not ( n74897 , n68838 );
buf ( n74898 , n74897 );
buf ( n74899 , n68634 );
or ( n74900 , n74509 , n74867 );
nand ( n74901 , n74867 , n69500 );
nand ( n74902 , n74900 , n74901 );
buf ( n74903 , n74902 );
buf ( n74904 , 1'b0 );
not ( n74905 , n68838 );
buf ( n8767 , n74905 );
buf ( n74907 , n68634 );
or ( n74908 , n74531 , n74867 );
nand ( n74909 , n74867 , n69477 );
nand ( n74910 , n74908 , n74909 );
buf ( n74911 , n74910 );
buf ( n74912 , 1'b0 );
not ( n74913 , n68838 );
buf ( n74914 , n74913 );
buf ( n74915 , n68634 );
not ( n74916 , n74551 );
or ( n74917 , n74916 , n74867 );
or ( n74918 , n74866 , n69448 );
nand ( n74919 , n74917 , n74918 );
buf ( n74920 , n74919 );
buf ( n74921 , 1'b0 );
not ( n74922 , n68838 );
buf ( n74923 , n74922 );
buf ( n8785 , n68634 );
and ( n74925 , n74867 , n3799 );
not ( n74926 , n74867 );
and ( n74927 , n74926 , n73928 );
or ( n74928 , n74925 , n74927 );
buf ( n74929 , n74928 );
buf ( n8791 , 1'b0 );
not ( n74931 , n68838 );
buf ( n8793 , n74931 );
buf ( n8794 , n68634 );
or ( n74934 , n74570 , n74867 );
or ( n74935 , n74866 , n69905 );
nand ( n74936 , n74934 , n74935 );
buf ( n8798 , n74936 );
buf ( n74938 , 1'b0 );
not ( n74939 , n68838 );
buf ( n74940 , n74939 );
buf ( n8802 , n68634 );
or ( n74942 , n74590 , n74867 );
nand ( n74943 , n74867 , n70063 );
nand ( n74944 , n74942 , n74943 );
buf ( n8806 , n74944 );
buf ( n8807 , 1'b0 );
not ( n74947 , n68838 );
buf ( n8809 , n74947 );
buf ( n74949 , n68634 );
or ( n74950 , n74612 , n74867 );
nand ( n74951 , n74867 , n69732 );
nand ( n74952 , n74950 , n74951 );
buf ( n8814 , n74952 );
buf ( n8815 , 1'b0 );
not ( n74955 , n68838 );
buf ( n74956 , n74955 );
buf ( n74957 , n68634 );
or ( n74958 , n74634 , n74867 );
nand ( n74959 , n74867 , n69725 );
nand ( n74960 , n74958 , n74959 );
buf ( n74961 , n74960 );
buf ( n74962 , 1'b0 );
not ( n74963 , n68838 );
buf ( n8825 , n74963 );
buf ( n74965 , n68634 );
not ( n74966 , n69697 );
and ( n74967 , n74867 , n74966 );
not ( n74968 , n74867 );
and ( n74969 , n74968 , n74654 );
nor ( n74970 , n74967 , n74969 );
buf ( n74971 , n74970 );
buf ( n74972 , 1'b0 );
not ( n74973 , n68838 );
buf ( n8835 , n74973 );
buf ( n8836 , n68634 );
or ( n74976 , n74674 , n74867 );
nand ( n74977 , n74867 , n69681 );
nand ( n74978 , n74976 , n74977 );
buf ( n8840 , n74978 );
buf ( n8841 , 1'b0 );
not ( n74981 , n68838 );
buf ( n74982 , n74981 );
buf ( n74983 , n68634 );
or ( n74984 , n74694 , n74867 );
nand ( n74985 , n74867 , n69842 );
nand ( n74986 , n74984 , n74985 );
buf ( n74987 , n74986 );
buf ( n74988 , 1'b0 );
not ( n74989 , n68838 );
buf ( n74990 , n74989 );
buf ( n74991 , n68634 );
or ( n74992 , n74714 , n74867 );
nand ( n74993 , n74867 , n69923 );
nand ( n74994 , n74992 , n74993 );
buf ( n74995 , n74994 );
buf ( n74996 , 1'b0 );
not ( n74997 , n68838 );
buf ( n8859 , n74997 );
buf ( n8860 , n68634 );
or ( n75000 , n74734 , n74867 );
nand ( n75001 , n74867 , n69761 );
nand ( n75002 , n75000 , n75001 );
buf ( n75003 , n75002 );
buf ( n8865 , 1'b0 );
not ( n75005 , n68838 );
buf ( n8867 , n75005 );
buf ( n8868 , n68634 );
or ( n75008 , n74754 , n74867 );
nand ( n75009 , n74867 , n69788 );
nand ( n75010 , n75008 , n75009 );
buf ( n8872 , n75010 );
buf ( n75012 , 1'b0 );
not ( n75013 , n68838 );
buf ( n75014 , n75013 );
buf ( n8876 , n68634 );
or ( n75016 , n74774 , n74867 );
nand ( n75017 , n74867 , n69892 );
nand ( n75018 , n75016 , n75017 );
buf ( n8880 , n75018 );
buf ( n8881 , 1'b0 );
not ( n75021 , n68838 );
buf ( n8883 , n75021 );
buf ( n75023 , n68634 );
or ( n75024 , n74796 , n74867 );
nand ( n75025 , n74867 , n69867 );
nand ( n75026 , n75024 , n75025 );
buf ( n8888 , n75026 );
buf ( n8889 , 1'b0 );
not ( n75029 , n68838 );
buf ( n75030 , n75029 );
buf ( n75031 , n68634 );
or ( n75032 , n74815 , n74867 );
nand ( n75033 , n74867 , n70045 );
nand ( n75034 , n75032 , n75033 );
buf ( n75035 , n75034 );
buf ( n75036 , 1'b0 );
not ( n75037 , n68838 );
buf ( n8899 , n75037 );
buf ( n75039 , n68634 );
or ( n75040 , n71207 , n74867 );
nand ( n75041 , n74867 , n69796 );
nand ( n75042 , n75040 , n75041 );
buf ( n8904 , n75042 );
buf ( n75044 , 1'b0 );
not ( n75045 , n68838 );
buf ( n75046 , n75045 );
buf ( n75047 , n68634 );
or ( n75048 , n71263 , n74867 );
nand ( n75049 , n74867 , n69815 );
nand ( n75050 , n75048 , n75049 );
buf ( n75051 , n75050 );
buf ( n75052 , 1'b0 );
not ( n75053 , n68838 );
buf ( n8915 , n75053 );
buf ( n75055 , n68634 );
or ( n75056 , n71319 , n74867 );
nand ( n75057 , n74867 , n69645 );
nand ( n75058 , n75056 , n75057 );
buf ( n75059 , n75058 );
buf ( n75060 , 1'b0 );
not ( n75061 , n68838 );
buf ( n75062 , n75061 );
buf ( n75063 , n68634 );
or ( n75064 , n71341 , n74867 );
nand ( n75065 , n74867 , n69630 );
nand ( n75066 , n75064 , n75065 );
buf ( n75067 , n75066 );
buf ( n75068 , 1'b0 );
not ( n75069 , n68838 );
buf ( n75070 , n75069 );
buf ( n75071 , n68634 );
or ( n75072 , n71435 , n74867 );
nand ( n75073 , n74867 , n69611 );
nand ( n75074 , n75072 , n75073 );
buf ( n75075 , n75074 );
buf ( n75076 , 1'b0 );
not ( n75077 , n68838 );
buf ( n8939 , n75077 );
buf ( n8940 , n68634 );
or ( n75080 , n71508 , n74867 );
nand ( n75081 , n74867 , n69597 );
nand ( n75082 , n75080 , n75081 );
buf ( n75083 , n75082 );
buf ( n8945 , 1'b0 );
not ( n75085 , n68838 );
buf ( n75086 , n75085 );
buf ( n75087 , n68634 );
or ( n75088 , n74836 , n74867 );
nand ( n75089 , n74867 , n69572 );
nand ( n75090 , n75088 , n75089 );
buf ( n75091 , n75090 );
buf ( n75092 , 1'b0 );
not ( n75093 , n68838 );
buf ( n8955 , n75093 );
buf ( n8956 , n68634 );
or ( n75096 , n71574 , n74867 );
nand ( n75097 , n74867 , n69585 );
nand ( n75098 , n75096 , n75097 );
buf ( n75099 , n75098 );
buf ( n8961 , 1'b0 );
not ( n75101 , n68838 );
buf ( n8963 , n75101 );
buf ( n8964 , n68634 );
or ( n75104 , n71654 , n74867 );
nand ( n75105 , n74867 , n69517 );
nand ( n75106 , n75104 , n75105 );
buf ( n75107 , n75106 );
buf ( n75108 , 1'b0 );
not ( n75109 , n68838 );
buf ( n75110 , n75109 );
buf ( n8972 , n68634 );
or ( n75112 , n71714 , n74867 );
nand ( n75113 , n74867 , n69529 );
nand ( n75114 , n75112 , n75113 );
buf ( n75115 , n75114 );
buf ( n8977 , 1'b0 );
not ( n75117 , n68838 );
buf ( n75118 , n75117 );
buf ( n75119 , n68634 );
or ( n75120 , n74856 , n74867 );
or ( n75121 , n74866 , n69962 );
nand ( n75122 , n75120 , n75121 );
buf ( n8984 , n75122 );
buf ( n75124 , 1'b0 );
not ( n75125 , n68838 );
buf ( n75126 , n75125 );
buf ( n8988 , n68634 );
and ( n75128 , n71843 , n2669 );
not ( n75129 , n71843 );
and ( n75130 , n75129 , n70082 );
or ( n75131 , n75128 , n75130 );
buf ( n75132 , n75131 );
buf ( n75133 , 1'b0 );
not ( n75134 , n68838 );
buf ( n75135 , n75134 );
buf ( n75136 , n68634 );
and ( n75137 , n71843 , n68810 );
not ( n75138 , n71843 );
and ( n75139 , n75138 , n70090 );
or ( n75140 , n75137 , n75139 );
buf ( n75141 , n75140 );
buf ( n75142 , 1'b0 );
not ( n75143 , n68838 );
buf ( n75144 , n75143 );
buf ( n75145 , n68634 );
and ( n75146 , n71843 , n2673 );
not ( n75147 , n71843 );
and ( n75148 , n75147 , n70031 );
or ( n75149 , n75146 , n75148 );
buf ( n75150 , n75149 );
buf ( n75151 , 1'b0 );
not ( n75152 , n68838 );
buf ( n9014 , n75152 );
buf ( n9015 , n68634 );
and ( n75155 , n71843 , n68814 );
not ( n75156 , n71843 );
and ( n75157 , n75156 , n70024 );
or ( n75158 , n75155 , n75157 );
buf ( n9020 , n75158 );
buf ( n75160 , 1'b0 );
not ( n75161 , n68838 );
buf ( n75162 , n75161 );
buf ( n9024 , n68634 );
and ( n75164 , n71725 , n68818 );
not ( n75165 , n71725 );
and ( n75166 , n75165 , n70038 );
or ( n75167 , n75164 , n75166 );
buf ( n9029 , n75167 );
buf ( n9030 , 1'b0 );
not ( n75170 , n68838 );
buf ( n75171 , n75170 );
buf ( n75172 , n68634 );
not ( n75173 , n71725 );
not ( n75174 , n75173 );
not ( n75175 , n70040 );
or ( n75176 , n75174 , n75175 );
nand ( n75177 , n71843 , n68823 );
nand ( n75178 , n75176 , n75177 );
buf ( n75179 , n75178 );
buf ( n75180 , 1'b0 );
not ( n75181 , n68838 );
buf ( n75182 , n75181 );
buf ( n75183 , n68634 );
and ( n75184 , n71725 , n68764 );
not ( n75185 , n71725 );
and ( n75186 , n75185 , n73902 );
or ( n75187 , n75184 , n75186 );
buf ( n75188 , n75187 );
buf ( n75189 , 1'b0 );
not ( n75190 , n68838 );
buf ( n9052 , n75190 );
buf ( n75192 , n68634 );
not ( n75193 , n70073 );
not ( n75194 , n71725 );
not ( n75195 , n75194 );
or ( n75196 , n75193 , n75195 );
not ( n75197 , n68826 );
or ( n75198 , n71842 , n75197 );
nand ( n75199 , n75196 , n75198 );
buf ( n75200 , n75199 );
buf ( n9062 , 1'b0 );
not ( n75202 , n68838 );
buf ( n75203 , n75202 );
buf ( n75204 , n68634 );
and ( n75205 , n71725 , n68766 );
not ( n75206 , n71725 );
and ( n75207 , n75206 , n72463 );
or ( n75208 , n75205 , n75207 );
buf ( n75209 , n75208 );
buf ( n75210 , 1'b0 );
not ( n75211 , n68838 );
buf ( n75212 , n75211 );
buf ( n75213 , n68634 );
and ( n75214 , n71725 , n2629 );
not ( n75215 , n71725 );
and ( n75216 , n75215 , n72452 );
or ( n75217 , n75214 , n75216 );
buf ( n75218 , n75217 );
buf ( n75219 , 1'b0 );
not ( n75220 , n68838 );
buf ( n9082 , n75220 );
buf ( n9083 , n68634 );
not ( n75223 , n70053 );
not ( n75224 , n75194 );
or ( n75225 , n75223 , n75224 );
not ( n75226 , n71725 );
not ( n75227 , n2689 );
or ( n75228 , n75226 , n75227 );
nand ( n75229 , n75225 , n75228 );
buf ( n9091 , n75229 );
buf ( n75231 , 1'b0 );
not ( n75232 , n68838 );
buf ( n75233 , n75232 );
buf ( n75234 , n68634 );
not ( n75235 , n69967 );
not ( n75236 , n71725 );
not ( n75237 , n75236 );
or ( n75238 , n75235 , n75237 );
not ( n75239 , n68830 );
or ( n75240 , n75226 , n75239 );
nand ( n75241 , n75238 , n75240 );
buf ( n75242 , n75241 );
buf ( n75243 , 1'b0 );
not ( n75244 , n68838 );
buf ( n75245 , n75244 );
buf ( n75246 , n68634 );
nor ( n75247 , n70861 , n70147 );
not ( n75248 , n75247 );
or ( n75249 , n75248 , n70181 );
or ( n75250 , n75247 , n70170 );
nand ( n75251 , n75249 , n75250 );
buf ( n75252 , n75251 );
buf ( n75253 , 1'b0 );
not ( n75254 , n68838 );
buf ( n75255 , n75254 );
buf ( n75256 , n68634 );
or ( n75257 , n75248 , n74865 );
not ( n75258 , n70161 );
or ( n75259 , n75247 , n75258 );
nand ( n75260 , n75257 , n75259 );
buf ( n75261 , n75260 );
buf ( n75262 , 1'b0 );
not ( n75263 , n68838 );
buf ( n9125 , n75263 );
buf ( n9126 , n68634 );
not ( n75266 , n70195 );
not ( n75267 , n70140 );
or ( n75268 , n75266 , n75267 );
nand ( n75269 , n70147 , n70139 );
nand ( n75270 , n75268 , n75269 );
not ( n75271 , n70217 );
and ( n75272 , n69358 , n75271 );
and ( n75273 , n75270 , n75272 );
nand ( n75274 , n75273 , n69123 );
and ( n75275 , n69357 , n75271 );
nand ( n75276 , n75270 , n75275 );
not ( n75277 , n75276 );
nor ( n75278 , n69123 , n69533 );
not ( n75279 , n75278 );
nand ( n75280 , n69123 , n69533 );
nand ( n75281 , n75279 , n75280 );
not ( n75282 , n75281 );
or ( n75283 , n3276 , n69059 );
not ( n75284 , n75283 );
not ( n75285 , n69010 );
not ( n75286 , n75285 );
nor ( n75287 , n75286 , n3320 );
nor ( n75288 , n75284 , n75287 );
not ( n75289 , n69025 );
not ( n75290 , n75289 );
nor ( n75291 , n75290 , n3350 );
nand ( n75292 , n69083 , n3346 );
or ( n75293 , n75291 , n75292 );
nand ( n75294 , n75290 , n3350 );
nand ( n75295 , n75293 , n75294 );
and ( n75296 , n75288 , n75295 );
nand ( n75297 , n69059 , n3276 );
or ( n75298 , n75287 , n75297 );
nand ( n75299 , n75286 , n3320 );
nand ( n75300 , n75298 , n75299 );
nor ( n75301 , n75296 , n75300 );
nor ( n75302 , n69083 , n3346 );
nor ( n75303 , n75291 , n75302 );
nor ( n75304 , n69072 , n69437 );
nand ( n75305 , n69095 , n70058 );
or ( n75306 , n75304 , n75305 );
nand ( n75307 , n69072 , n69437 );
nand ( n75308 , n75306 , n75307 );
or ( n75309 , n70058 , n69095 );
and ( n75310 , n3815 , n2728 );
xor ( n75311 , n70051 , n75310 );
and ( n75312 , n75311 , n69106 );
and ( n75313 , n70051 , n75310 );
or ( n75314 , n75312 , n75313 );
nand ( n75315 , n75309 , n75314 );
nor ( n75316 , n75304 , n75315 );
or ( n75317 , n75308 , n75316 );
nand ( n75318 , n75288 , n75303 , n75317 );
nand ( n75319 , n75301 , n75318 );
not ( n75320 , n75319 );
nor ( n75321 , n68988 , n3405 );
or ( n75322 , n75320 , n75321 );
nand ( n75323 , n68988 , n3405 );
nand ( n75324 , n75322 , n75323 );
not ( n75325 , n75324 );
or ( n75326 , n75282 , n75325 );
or ( n75327 , n75324 , n75281 );
nand ( n75328 , n75326 , n75327 );
nand ( n75329 , n75277 , n75328 );
not ( n75330 , n69357 );
nor ( n75331 , n75330 , n75271 );
and ( n75332 , n75270 , n75331 );
nor ( n75333 , n69123 , n69535 );
not ( n75334 , n75333 );
nand ( n75335 , n69123 , n69535 );
nand ( n75336 , n75334 , n75335 );
not ( n75337 , n75336 );
or ( n75338 , n3282 , n69059 );
not ( n75339 , n75338 );
not ( n75340 , n75285 );
nor ( n75341 , n75340 , n3316 );
nor ( n75342 , n75339 , n75341 );
not ( n75343 , n75289 );
nor ( n75344 , n75343 , n69492 );
nand ( n75345 , n69083 , n3342 );
or ( n75346 , n75344 , n75345 );
nand ( n75347 , n75343 , n69492 );
nand ( n75348 , n75346 , n75347 );
and ( n75349 , n75342 , n75348 );
nand ( n75350 , n69059 , n3282 );
or ( n75351 , n75341 , n75350 );
nand ( n75352 , n75340 , n3316 );
nand ( n75353 , n75351 , n75352 );
nor ( n75354 , n75349 , n75353 );
nor ( n75355 , n69083 , n3342 );
nor ( n75356 , n75344 , n75355 );
nor ( n75357 , n69072 , n3301 );
nand ( n75358 , n69095 , n70069 );
or ( n75359 , n75357 , n75358 );
nand ( n75360 , n69072 , n3301 );
nand ( n75361 , n75359 , n75360 );
or ( n75362 , n70069 , n69095 );
and ( n75363 , n69957 , n2728 );
xor ( n75364 , n70049 , n75363 );
and ( n75365 , n75364 , n69106 );
and ( n75366 , n70049 , n75363 );
or ( n75367 , n75365 , n75366 );
nand ( n75368 , n75362 , n75367 );
nor ( n75369 , n75357 , n75368 );
or ( n75370 , n75361 , n75369 );
nand ( n75371 , n75342 , n75356 , n75370 );
nand ( n75372 , n75354 , n75371 );
not ( n75373 , n75372 );
nor ( n75374 , n68988 , n69546 );
or ( n75375 , n75373 , n75374 );
nand ( n75376 , n68988 , n69546 );
nand ( n75377 , n75375 , n75376 );
not ( n75378 , n75377 );
or ( n75379 , n75337 , n75378 );
or ( n75380 , n75377 , n75336 );
nand ( n75381 , n75379 , n75380 );
nand ( n75382 , n75332 , n75381 );
nor ( n75383 , n70136 , n70147 );
not ( n75384 , n70195 );
and ( n75385 , n75384 , n70863 );
nor ( n75386 , n69357 , n75271 );
nor ( n75387 , n75385 , n75386 );
or ( n75388 , n75383 , n75387 , n71992 );
not ( n75389 , n75388 );
and ( n75390 , n75389 , n68720 );
not ( n75391 , n72020 );
nor ( n75392 , n75390 , n75391 );
nand ( n75393 , n75274 , n75329 , n75382 , n75392 );
buf ( n75394 , n75393 );
buf ( n9256 , 1'b0 );
not ( n75396 , n68838 );
buf ( n9258 , n75396 );
buf ( n9259 , n68634 );
nand ( n75399 , n75273 , n68988 );
not ( n75400 , n75321 );
nand ( n75401 , n75400 , n75323 );
not ( n75402 , n75401 );
not ( n75403 , n75319 );
or ( n75404 , n75402 , n75403 );
or ( n75405 , n75319 , n75401 );
nand ( n75406 , n75404 , n75405 );
nand ( n75407 , n75277 , n75406 );
not ( n75408 , n75374 );
nand ( n75409 , n75408 , n75376 );
not ( n75410 , n75409 );
not ( n75411 , n75372 );
or ( n75412 , n75410 , n75411 );
or ( n75413 , n75372 , n75409 );
nand ( n75414 , n75412 , n75413 );
nand ( n75415 , n75332 , n75414 );
and ( n75416 , n75389 , n68725 );
nor ( n75417 , n75416 , n72072 );
nand ( n75418 , n75399 , n75407 , n75415 , n75417 );
buf ( n75419 , n75418 );
buf ( n75420 , 1'b0 );
not ( n75421 , n68838 );
buf ( n9283 , n75421 );
buf ( n9284 , n68634 );
nand ( n75424 , n75273 , n69010 );
not ( n75425 , n75299 );
nor ( n75426 , n75425 , n75287 );
not ( n75427 , n75426 );
and ( n75428 , n75303 , n75317 , n75283 );
not ( n75429 , n75283 );
not ( n75430 , n75295 );
or ( n75431 , n75429 , n75430 );
nand ( n75432 , n75431 , n75297 );
nor ( n75433 , n75428 , n75432 );
not ( n75434 , n75433 );
or ( n75435 , n75427 , n75434 );
or ( n75436 , n75433 , n75426 );
nand ( n75437 , n75435 , n75436 );
nand ( n75438 , n75277 , n75437 );
not ( n75439 , n75352 );
nor ( n75440 , n75439 , n75341 );
not ( n75441 , n75440 );
and ( n75442 , n75356 , n75370 , n75338 );
not ( n75443 , n75338 );
not ( n75444 , n75348 );
or ( n75445 , n75443 , n75444 );
nand ( n75446 , n75445 , n75350 );
nor ( n75447 , n75442 , n75446 );
not ( n75448 , n75447 );
or ( n75449 , n75441 , n75448 );
or ( n75450 , n75447 , n75440 );
nand ( n75451 , n75449 , n75450 );
nand ( n75452 , n75332 , n75451 );
and ( n75453 , n75389 , n68730 );
nor ( n75454 , n75453 , n72138 );
nand ( n75455 , n75424 , n75438 , n75452 , n75454 );
buf ( n9317 , n75455 );
buf ( n9318 , 1'b0 );
not ( n75458 , n68838 );
buf ( n75459 , n75458 );
buf ( n75460 , n68634 );
nand ( n75461 , n75273 , n69059 );
and ( n75462 , n75283 , n75297 );
not ( n75463 , n75462 );
and ( n75464 , n75303 , n75317 );
nor ( n75465 , n75464 , n75295 );
not ( n75466 , n75465 );
or ( n75467 , n75463 , n75466 );
or ( n75468 , n75465 , n75462 );
nand ( n75469 , n75467 , n75468 );
nand ( n75470 , n75277 , n75469 );
and ( n75471 , n75338 , n75350 );
not ( n75472 , n75471 );
and ( n75473 , n75356 , n75370 );
nor ( n75474 , n75473 , n75348 );
not ( n75475 , n75474 );
or ( n75476 , n75472 , n75475 );
or ( n75477 , n75474 , n75471 );
nand ( n75478 , n75476 , n75477 );
nand ( n75479 , n75332 , n75478 );
and ( n75480 , n75389 , n68735 );
nor ( n75481 , n75480 , n72200 );
nand ( n75482 , n75461 , n75470 , n75479 , n75481 );
buf ( n75483 , n75482 );
buf ( n75484 , 1'b0 );
not ( n75485 , n68838 );
buf ( n75486 , n75485 );
buf ( n75487 , n68634 );
nand ( n75488 , n75273 , n69025 );
not ( n75489 , n75291 );
nand ( n75490 , n75489 , n75294 );
not ( n75491 , n75490 );
not ( n75492 , n75317 );
or ( n75493 , n75492 , n75302 );
nand ( n75494 , n75493 , n75292 );
not ( n75495 , n75494 );
or ( n75496 , n75491 , n75495 );
or ( n75497 , n75494 , n75490 );
nand ( n75498 , n75496 , n75497 );
nand ( n75499 , n75277 , n75498 );
not ( n75500 , n75344 );
nand ( n75501 , n75500 , n75347 );
not ( n75502 , n75501 );
not ( n75503 , n75370 );
or ( n75504 , n75503 , n75355 );
nand ( n75505 , n75504 , n75345 );
not ( n75506 , n75505 );
or ( n75507 , n75502 , n75506 );
or ( n75508 , n75505 , n75501 );
nand ( n75509 , n75507 , n75508 );
nand ( n75510 , n75332 , n75509 );
and ( n75511 , n75389 , n68740 );
nor ( n75512 , n75511 , n72262 );
nand ( n75513 , n75488 , n75499 , n75510 , n75512 );
buf ( n75514 , n75513 );
buf ( n75515 , 1'b0 );
not ( n75516 , n68838 );
buf ( n75517 , n75516 );
buf ( n75518 , n68634 );
nand ( n75519 , n75273 , n69083 );
not ( n75520 , n75292 );
nor ( n75521 , n75520 , n75302 );
not ( n75522 , n75521 );
not ( n75523 , n75492 );
or ( n75524 , n75522 , n75523 );
or ( n75525 , n75492 , n75521 );
nand ( n75526 , n75524 , n75525 );
nand ( n75527 , n75277 , n75526 );
not ( n75528 , n75345 );
nor ( n75529 , n75528 , n75355 );
not ( n75530 , n75529 );
not ( n75531 , n75503 );
or ( n75532 , n75530 , n75531 );
or ( n75533 , n75503 , n75529 );
nand ( n75534 , n75532 , n75533 );
nand ( n75535 , n75332 , n75534 );
not ( n75536 , n75388 );
not ( n75537 , n2604 );
not ( n75538 , n75537 );
and ( n75539 , n75536 , n75538 );
not ( n75540 , n3815 );
not ( n75541 , n75275 );
or ( n75542 , n75540 , n75541 );
nand ( n75543 , n75331 , n69957 );
nand ( n75544 , n75542 , n75543 );
xnor ( n75545 , n75544 , n2728 );
or ( n75546 , n71725 , n75545 );
nand ( n75547 , n75546 , n72311 );
nor ( n75548 , n75539 , n75547 );
nand ( n75549 , n75519 , n75527 , n75535 , n75548 );
buf ( n75550 , n75549 );
buf ( n75551 , 1'b0 );
not ( n75552 , n68838 );
buf ( n75553 , n75552 );
buf ( n9415 , n68634 );
nand ( n75555 , n75273 , n69072 );
nand ( n75556 , n75315 , n75305 );
not ( n75557 , n75556 );
not ( n75558 , n75304 );
nand ( n75559 , n75558 , n75307 );
not ( n75560 , n75559 );
or ( n75561 , n75557 , n75560 );
or ( n75562 , n75559 , n75556 );
nand ( n75563 , n75561 , n75562 );
nand ( n75564 , n75277 , n75563 );
nand ( n75565 , n75368 , n75358 );
not ( n75566 , n75565 );
not ( n75567 , n75357 );
nand ( n75568 , n75567 , n75360 );
not ( n75569 , n75568 );
or ( n75570 , n75566 , n75569 );
or ( n75571 , n75568 , n75565 );
nand ( n75572 , n75570 , n75571 );
nand ( n75573 , n75332 , n75572 );
and ( n75574 , n75389 , n68747 );
nor ( n75575 , n75574 , n72368 );
nand ( n75576 , n75555 , n75564 , n75573 , n75575 );
buf ( n75577 , n75576 );
buf ( n75578 , 1'b0 );
not ( n75579 , n68838 );
buf ( n75580 , n75579 );
buf ( n75581 , n68634 );
not ( n75582 , n75314 );
nand ( n75583 , n75305 , n75309 );
not ( n75584 , n75583 );
or ( n75585 , n75582 , n75584 );
or ( n75586 , n75583 , n75314 );
nand ( n75587 , n75585 , n75586 );
nand ( n75588 , n75277 , n75587 );
nand ( n75589 , n75273 , n69095 );
not ( n75590 , n75367 );
nand ( n75591 , n75358 , n75362 );
not ( n75592 , n75591 );
or ( n75593 , n75590 , n75592 );
or ( n75594 , n75591 , n75367 );
nand ( n75595 , n75593 , n75594 );
nand ( n75596 , n75332 , n75595 );
not ( n75597 , n75388 );
not ( n75598 , n68750 );
not ( n75599 , n75598 );
and ( n75600 , n75597 , n75599 );
not ( n75601 , n70859 );
not ( n75602 , n3915 );
or ( n75603 , n75601 , n75602 );
nand ( n75604 , n75603 , n75546 );
nor ( n75605 , n75600 , n75604 );
nand ( n75606 , n75588 , n75589 , n75596 , n75605 );
buf ( n75607 , n75606 );
buf ( n75608 , 1'b0 );
not ( n75609 , n68838 );
buf ( n75610 , n75609 );
buf ( n75611 , n68634 );
nand ( n75612 , n75273 , n69106 );
xor ( n75613 , n70051 , n75310 );
xor ( n75614 , n75613 , n69106 );
nand ( n75615 , n75277 , n75614 );
xor ( n75616 , n70049 , n75363 );
xor ( n75617 , n75616 , n69106 );
nand ( n75618 , n75332 , n75617 );
and ( n75619 , n75389 , n68754 );
and ( n75620 , n70041 , n70859 );
nor ( n75621 , n75619 , n75620 );
nand ( n75622 , n75612 , n75615 , n75618 , n75621 );
buf ( n75623 , n75622 );
buf ( n75624 , 1'b0 );
not ( n75625 , n68838 );
buf ( n9487 , n75625 );
buf ( n9488 , n68634 );
nand ( n75628 , n75273 , n69240 );
not ( n75629 , n69240 );
not ( n75630 , n69798 );
and ( n75631 , n75629 , n75630 );
and ( n75632 , n69240 , n69798 );
nor ( n75633 , n75631 , n75632 );
not ( n75634 , n75633 );
or ( n75635 , n69045 , n69522 );
not ( n75636 , n75635 );
nor ( n75637 , n68977 , n69507 );
nor ( n75638 , n75636 , n75637 );
or ( n75639 , n75278 , n75323 );
nand ( n75640 , n75639 , n75280 );
and ( n75641 , n75638 , n75640 );
nand ( n75642 , n69045 , n69522 );
or ( n75643 , n75637 , n75642 );
nand ( n75644 , n68977 , n69507 );
nand ( n75645 , n75643 , n75644 );
nor ( n75646 , n75641 , n75645 );
nor ( n75647 , n75278 , n75321 );
and ( n75648 , n75638 , n75647 );
nand ( n75649 , n75648 , n75319 );
nand ( n75650 , n75646 , n75649 );
nor ( n75651 , n68934 , n3466 );
nor ( n75652 , n68961 , n3450 );
nor ( n75653 , n75651 , n75652 );
nor ( n75654 , n68947 , n69558 );
nor ( n75655 , n68908 , n69577 );
nor ( n75656 , n75654 , n75655 );
nand ( n75657 , n75653 , n75656 );
not ( n75658 , n75657 );
nor ( n75659 , n69157 , n69806 );
not ( n75660 , n75659 );
nor ( n75661 , n69176 , n69651 );
nor ( n75662 , n69187 , n2697 );
nor ( n75663 , n75661 , n75662 );
nand ( n75664 , n75660 , n75663 );
not ( n75665 , n75664 );
and ( n75666 , n75650 , n75658 , n75665 );
nand ( n75667 , n68908 , n69577 );
or ( n75668 , n75654 , n75667 );
nand ( n75669 , n68947 , n69558 );
nand ( n75670 , n75668 , n75669 );
and ( n75671 , n75653 , n75670 );
nand ( n75672 , n68961 , n3450 );
or ( n75673 , n75651 , n75672 );
nand ( n75674 , n68934 , n3466 );
nand ( n75675 , n75673 , n75674 );
nor ( n75676 , n75671 , n75675 );
or ( n75677 , n75676 , n75664 );
nand ( n75678 , n69187 , n2697 );
or ( n75679 , n75661 , n75678 );
nand ( n75680 , n69176 , n69651 );
nand ( n75681 , n75679 , n75680 );
not ( n75682 , n75681 );
or ( n75683 , n75659 , n75682 );
nand ( n75684 , n69157 , n69806 );
nand ( n75685 , n75677 , n75683 , n75684 );
nor ( n75686 , n75666 , n75685 );
not ( n75687 , n75686 );
or ( n75688 , n75634 , n75687 );
or ( n75689 , n75686 , n75633 );
nand ( n75690 , n75688 , n75689 );
nand ( n75691 , n75277 , n75690 );
not ( n75692 , n69240 );
not ( n75693 , n69800 );
and ( n75694 , n75692 , n75693 );
and ( n75695 , n69240 , n69800 );
nor ( n75696 , n75694 , n75695 );
not ( n75697 , n75696 );
or ( n75698 , n69045 , n69524 );
not ( n75699 , n75698 );
nor ( n75700 , n68977 , n69509 );
nor ( n75701 , n75699 , n75700 );
or ( n75702 , n75333 , n75376 );
nand ( n75703 , n75702 , n75335 );
and ( n75704 , n75701 , n75703 );
nand ( n75705 , n69045 , n69524 );
or ( n75706 , n75700 , n75705 );
nand ( n75707 , n68977 , n69509 );
nand ( n75708 , n75706 , n75707 );
nor ( n75709 , n75704 , n75708 );
nor ( n75710 , n75333 , n75374 );
and ( n75711 , n75701 , n75710 );
nand ( n75712 , n75711 , n75372 );
nand ( n75713 , n75709 , n75712 );
nor ( n75714 , n68934 , n69607 );
nor ( n75715 , n68961 , n69591 );
nor ( n75716 , n75714 , n75715 );
nor ( n75717 , n68947 , n69562 );
nor ( n75718 , n68908 , n69579 );
nor ( n75719 , n75717 , n75718 );
nand ( n75720 , n75716 , n75719 );
not ( n75721 , n75720 );
nor ( n75722 , n69157 , n69810 );
not ( n75723 , n75722 );
nor ( n75724 , n69176 , n3510 );
nor ( n75725 , n69187 , n3498 );
nor ( n75726 , n75724 , n75725 );
nand ( n75727 , n75723 , n75726 );
not ( n75728 , n75727 );
and ( n75729 , n75713 , n75721 , n75728 );
nand ( n75730 , n68908 , n69579 );
or ( n75731 , n75717 , n75730 );
nand ( n75732 , n68947 , n69562 );
nand ( n75733 , n75731 , n75732 );
and ( n75734 , n75716 , n75733 );
nand ( n75735 , n68961 , n69591 );
or ( n75736 , n75714 , n75735 );
nand ( n75737 , n68934 , n69607 );
nand ( n75738 , n75736 , n75737 );
nor ( n75739 , n75734 , n75738 );
or ( n75740 , n75739 , n75727 );
nand ( n75741 , n69187 , n3498 );
or ( n75742 , n75724 , n75741 );
nand ( n75743 , n69176 , n3510 );
nand ( n75744 , n75742 , n75743 );
not ( n75745 , n75744 );
or ( n75746 , n75722 , n75745 );
nand ( n75747 , n69157 , n69810 );
nand ( n75748 , n75740 , n75746 , n75747 );
nor ( n75749 , n75729 , n75748 );
not ( n75750 , n75749 );
or ( n75751 , n75697 , n75750 );
or ( n75752 , n75749 , n75696 );
nand ( n75753 , n75751 , n75752 );
nand ( n75754 , n75332 , n75753 );
and ( n75755 , n75389 , n68670 );
nor ( n75756 , n75755 , n73456 );
nand ( n75757 , n75628 , n75691 , n75754 , n75756 );
buf ( n9619 , n75757 );
buf ( n9620 , 1'b0 );
not ( n75760 , n68838 );
buf ( n9622 , n75760 );
buf ( n9623 , n68634 );
nand ( n75763 , n75273 , n69157 );
not ( n75764 , n75684 );
nor ( n75765 , n75764 , n75659 );
not ( n75766 , n75765 );
and ( n75767 , n75650 , n75658 , n75663 );
not ( n75768 , n75681 );
not ( n75769 , n75676 );
nand ( n75770 , n75769 , n75663 );
nand ( n75771 , n75768 , n75770 );
nor ( n75772 , n75767 , n75771 );
not ( n75773 , n75772 );
or ( n75774 , n75766 , n75773 );
or ( n75775 , n75772 , n75765 );
nand ( n75776 , n75774 , n75775 );
nand ( n75777 , n75277 , n75776 );
not ( n75778 , n75747 );
nor ( n75779 , n75778 , n75722 );
not ( n75780 , n75779 );
and ( n75781 , n75713 , n75721 , n75726 );
not ( n75782 , n75744 );
not ( n75783 , n75739 );
nand ( n75784 , n75783 , n75726 );
nand ( n75785 , n75782 , n75784 );
nor ( n75786 , n75781 , n75785 );
not ( n75787 , n75786 );
or ( n75788 , n75780 , n75787 );
or ( n75789 , n75786 , n75779 );
nand ( n75790 , n75788 , n75789 );
nand ( n75791 , n75332 , n75790 );
and ( n75792 , n75389 , n68675 );
nor ( n75793 , n75792 , n73478 );
nand ( n75794 , n75763 , n75777 , n75791 , n75793 );
buf ( n9656 , n75794 );
buf ( n75796 , 1'b0 );
not ( n75797 , n68838 );
buf ( n75798 , n75797 );
buf ( n75799 , n68634 );
nand ( n75800 , n75273 , n69176 );
not ( n75801 , n75661 );
nand ( n75802 , n75801 , n75680 );
not ( n75803 , n75802 );
or ( n75804 , n75676 , n75662 );
not ( n75805 , n75662 );
nand ( n75806 , n75805 , n75650 , n75658 );
nand ( n75807 , n75804 , n75806 , n75678 );
not ( n75808 , n75807 );
or ( n75809 , n75803 , n75808 );
or ( n75810 , n75807 , n75802 );
nand ( n75811 , n75809 , n75810 );
nand ( n75812 , n75277 , n75811 );
not ( n75813 , n75724 );
nand ( n75814 , n75813 , n75743 );
not ( n75815 , n75814 );
or ( n75816 , n75739 , n75725 );
not ( n75817 , n75725 );
nand ( n75818 , n75817 , n75713 , n75721 );
nand ( n75819 , n75816 , n75818 , n75741 );
not ( n75820 , n75819 );
or ( n75821 , n75815 , n75820 );
or ( n75822 , n75819 , n75814 );
nand ( n75823 , n75821 , n75822 );
nand ( n75824 , n75332 , n75823 );
and ( n75825 , n75389 , n68680 );
nor ( n75826 , n75825 , n73500 );
nand ( n75827 , n75800 , n75812 , n75824 , n75826 );
buf ( n9689 , n75827 );
buf ( n75829 , 1'b0 );
not ( n75830 , n68838 );
buf ( n75831 , n75830 );
buf ( n75832 , n68634 );
nand ( n75833 , n75273 , n69187 );
not ( n75834 , n75662 );
nand ( n75835 , n75834 , n75678 );
not ( n75836 , n75835 );
or ( n75837 , n75649 , n75657 );
or ( n75838 , n75657 , n75646 );
nand ( n75839 , n75837 , n75838 , n75676 );
not ( n75840 , n75839 );
or ( n75841 , n75836 , n75840 );
or ( n75842 , n75839 , n75835 );
nand ( n75843 , n75841 , n75842 );
nand ( n75844 , n75277 , n75843 );
not ( n75845 , n75725 );
nand ( n75846 , n75845 , n75741 );
not ( n75847 , n75846 );
or ( n75848 , n75712 , n75720 );
or ( n75849 , n75720 , n75709 );
nand ( n75850 , n75848 , n75849 , n75739 );
not ( n75851 , n75850 );
or ( n75852 , n75847 , n75851 );
or ( n75853 , n75850 , n75846 );
nand ( n75854 , n75852 , n75853 );
nand ( n75855 , n75332 , n75854 );
and ( n75856 , n75389 , n68685 );
nor ( n75857 , n75856 , n73521 );
nand ( n75858 , n75833 , n75844 , n75855 , n75857 );
buf ( n9720 , n75858 );
buf ( n9721 , 1'b0 );
not ( n75861 , n68838 );
buf ( n75862 , n75861 );
buf ( n75863 , n68634 );
nand ( n75864 , n75273 , n68934 );
not ( n75865 , n75674 );
nor ( n75866 , n75865 , n75651 );
not ( n75867 , n75866 );
not ( n75868 , n75652 );
and ( n75869 , n75656 , n75868 );
and ( n75870 , n75648 , n75869 , n75319 );
not ( n75871 , n75869 );
not ( n75872 , n75646 );
not ( n75873 , n75872 );
or ( n75874 , n75871 , n75873 );
and ( n75875 , n75670 , n75868 );
not ( n75876 , n75672 );
nor ( n75877 , n75875 , n75876 );
nand ( n75878 , n75874 , n75877 );
nor ( n75879 , n75870 , n75878 );
not ( n75880 , n75879 );
or ( n75881 , n75867 , n75880 );
or ( n75882 , n75879 , n75866 );
nand ( n75883 , n75881 , n75882 );
nand ( n75884 , n75277 , n75883 );
not ( n75885 , n75737 );
nor ( n75886 , n75885 , n75714 );
not ( n75887 , n75886 );
not ( n75888 , n75715 );
and ( n75889 , n75719 , n75888 );
and ( n75890 , n75711 , n75889 , n75372 );
not ( n75891 , n75889 );
not ( n75892 , n75709 );
not ( n75893 , n75892 );
or ( n75894 , n75891 , n75893 );
and ( n75895 , n75733 , n75888 );
not ( n75896 , n75735 );
nor ( n75897 , n75895 , n75896 );
nand ( n75898 , n75894 , n75897 );
nor ( n75899 , n75890 , n75898 );
not ( n75900 , n75899 );
or ( n75901 , n75887 , n75900 );
or ( n75902 , n75899 , n75886 );
nand ( n75903 , n75901 , n75902 );
nand ( n75904 , n75332 , n75903 );
and ( n75905 , n75389 , n68690 );
not ( n75906 , n73547 );
nor ( n75907 , n75905 , n75906 );
nand ( n75908 , n75864 , n75884 , n75904 , n75907 );
buf ( n75909 , n75908 );
buf ( n75910 , 1'b0 );
not ( n75911 , n68838 );
buf ( n75912 , n75911 );
buf ( n75913 , n68634 );
nand ( n75914 , n75273 , n68961 );
and ( n75915 , n75868 , n75672 );
not ( n75916 , n75915 );
and ( n75917 , n75872 , n75656 );
and ( n75918 , n75648 , n75319 , n75656 );
nor ( n75919 , n75917 , n75918 , n75670 );
not ( n75920 , n75919 );
or ( n75921 , n75916 , n75920 );
or ( n75922 , n75919 , n75915 );
nand ( n75923 , n75921 , n75922 );
nand ( n75924 , n75277 , n75923 );
and ( n75925 , n75888 , n75735 );
not ( n75926 , n75925 );
and ( n75927 , n75892 , n75719 );
and ( n75928 , n75711 , n75372 , n75719 );
nor ( n75929 , n75927 , n75928 , n75733 );
not ( n75930 , n75929 );
or ( n75931 , n75926 , n75930 );
or ( n75932 , n75929 , n75925 );
nand ( n75933 , n75931 , n75932 );
nand ( n75934 , n75332 , n75933 );
and ( n75935 , n75389 , n68695 );
not ( n75936 , n73571 );
nor ( n75937 , n75935 , n75936 );
nand ( n75938 , n75914 , n75924 , n75934 , n75937 );
buf ( n75939 , n75938 );
buf ( n75940 , 1'b0 );
not ( n75941 , n68838 );
buf ( n75942 , n75941 );
buf ( n75943 , n68634 );
nand ( n75944 , n75273 , n68947 );
not ( n75945 , n75654 );
nand ( n75946 , n75945 , n75669 );
not ( n75947 , n75946 );
or ( n75948 , n75646 , n75655 );
not ( n75949 , n75655 );
nand ( n75950 , n75949 , n75648 , n75319 );
nand ( n75951 , n75948 , n75950 , n75667 );
not ( n75952 , n75951 );
or ( n75953 , n75947 , n75952 );
or ( n75954 , n75951 , n75946 );
nand ( n75955 , n75953 , n75954 );
nand ( n75956 , n75277 , n75955 );
not ( n75957 , n75717 );
nand ( n75958 , n75957 , n75732 );
not ( n75959 , n75958 );
or ( n75960 , n75709 , n75718 );
not ( n75961 , n75718 );
nand ( n75962 , n75961 , n75711 , n75372 );
nand ( n75963 , n75960 , n75962 , n75730 );
not ( n75964 , n75963 );
or ( n75965 , n75959 , n75964 );
or ( n75966 , n75963 , n75958 );
nand ( n75967 , n75965 , n75966 );
nand ( n75968 , n75332 , n75967 );
and ( n75969 , n75389 , n68700 );
not ( n75970 , n73645 );
nor ( n75971 , n75969 , n75970 );
nand ( n75972 , n75944 , n75956 , n75968 , n75971 );
buf ( n75973 , n75972 );
buf ( n75974 , 1'b0 );
not ( n75975 , n68838 );
buf ( n75976 , n75975 );
buf ( n75977 , n68634 );
nand ( n75978 , n75273 , n68908 );
not ( n75979 , n75655 );
nand ( n75980 , n75979 , n75667 );
not ( n75981 , n75980 );
not ( n75982 , n75650 );
or ( n75983 , n75981 , n75982 );
or ( n75984 , n75650 , n75980 );
nand ( n75985 , n75983 , n75984 );
nand ( n75986 , n75277 , n75985 );
not ( n75987 , n75718 );
nand ( n75988 , n75987 , n75730 );
not ( n75989 , n75988 );
not ( n75990 , n75713 );
or ( n75991 , n75989 , n75990 );
or ( n75992 , n75713 , n75988 );
nand ( n75993 , n75991 , n75992 );
nand ( n75994 , n75332 , n75993 );
and ( n75995 , n75389 , n68705 );
not ( n75996 , n73670 );
nor ( n75997 , n75995 , n75996 );
nand ( n75998 , n75978 , n75986 , n75994 , n75997 );
buf ( n75999 , n75998 );
buf ( n76000 , 1'b0 );
not ( n76001 , n68838 );
buf ( n76002 , n76001 );
buf ( n76003 , n68634 );
nand ( n76004 , n75273 , n68977 );
not ( n76005 , n75644 );
nor ( n76006 , n76005 , n75637 );
not ( n76007 , n76006 );
and ( n76008 , n75319 , n75647 , n75635 );
not ( n76009 , n75635 );
not ( n76010 , n75640 );
or ( n76011 , n76009 , n76010 );
nand ( n76012 , n76011 , n75642 );
nor ( n76013 , n76008 , n76012 );
not ( n76014 , n76013 );
or ( n76015 , n76007 , n76014 );
or ( n76016 , n76013 , n76006 );
nand ( n76017 , n76015 , n76016 );
nand ( n76018 , n75277 , n76017 );
not ( n76019 , n75707 );
nor ( n76020 , n76019 , n75700 );
not ( n76021 , n76020 );
and ( n76022 , n75372 , n75710 , n75698 );
not ( n76023 , n75698 );
not ( n76024 , n75703 );
or ( n76025 , n76023 , n76024 );
nand ( n76026 , n76025 , n75705 );
nor ( n76027 , n76022 , n76026 );
not ( n76028 , n76027 );
or ( n76029 , n76021 , n76028 );
or ( n76030 , n76027 , n76020 );
nand ( n76031 , n76029 , n76030 );
nand ( n76032 , n75332 , n76031 );
and ( n76033 , n75389 , n68710 );
not ( n76034 , n73694 );
nor ( n76035 , n76033 , n76034 );
nand ( n76036 , n76004 , n76018 , n76032 , n76035 );
buf ( n76037 , n76036 );
buf ( n76038 , 1'b0 );
not ( n76039 , n68838 );
buf ( n76040 , n76039 );
buf ( n76041 , n68634 );
nand ( n76042 , n75273 , n69045 );
and ( n76043 , n75635 , n75642 );
not ( n76044 , n76043 );
and ( n76045 , n75319 , n75647 );
nor ( n76046 , n76045 , n75640 );
not ( n76047 , n76046 );
or ( n76048 , n76044 , n76047 );
or ( n76049 , n76046 , n76043 );
nand ( n76050 , n76048 , n76049 );
nand ( n76051 , n75277 , n76050 );
and ( n76052 , n75698 , n75705 );
not ( n76053 , n76052 );
and ( n76054 , n75372 , n75710 );
nor ( n76055 , n76054 , n75703 );
not ( n76056 , n76055 );
or ( n76057 , n76053 , n76056 );
or ( n76058 , n76055 , n76052 );
nand ( n76059 , n76057 , n76058 );
nand ( n76060 , n75332 , n76059 );
and ( n76061 , n75389 , n68715 );
not ( n76062 , n73719 );
nor ( n76063 , n76061 , n76062 );
nand ( n76064 , n76042 , n76051 , n76060 , n76063 );
buf ( n76065 , n76064 );
buf ( n76066 , 1'b0 );
not ( n76067 , n68838 );
buf ( n76068 , n76067 );
buf ( n76069 , n68634 );
nand ( n76070 , n75273 , n2728 );
xor ( n76071 , n3815 , n2728 );
nand ( n76072 , n75277 , n76071 );
xor ( n76073 , n69957 , n2728 );
nand ( n76074 , n75332 , n76073 );
and ( n76075 , n75389 , n68759 );
and ( n76076 , n69950 , n70859 );
nor ( n76077 , n76075 , n76076 );
nand ( n76078 , n76070 , n76072 , n76074 , n76077 );
buf ( n76079 , n76078 );
buf ( n76080 , 1'b0 );
not ( n76081 , n68838 );
buf ( n9943 , n76081 );
buf ( n9944 , n68634 );
not ( n76084 , n69123 );
or ( n76085 , n71992 , n76084 );
nand ( n76086 , n70859 , n2519 );
nand ( n76087 , n76085 , n76086 );
buf ( n9949 , n76087 );
buf ( n9950 , 1'b0 );
not ( n76090 , n68838 );
buf ( n9952 , n76090 );
buf ( n9953 , n68634 );
not ( n76093 , n68988 );
or ( n76094 , n71992 , n76093 );
not ( n76095 , n68659 );
or ( n76096 , n72071 , n76095 );
nand ( n76097 , n76094 , n76096 );
buf ( n76098 , n76097 );
buf ( n76099 , 1'b0 );
not ( n76100 , n68838 );
buf ( n76101 , n76100 );
buf ( n76102 , n68634 );
not ( n76103 , n69010 );
not ( n76104 , n70139 );
or ( n76105 , n76103 , n76104 );
nand ( n76106 , n70859 , n68660 );
nand ( n76107 , n76105 , n76106 );
buf ( n76108 , n76107 );
buf ( n76109 , 1'b0 );
not ( n76110 , n68838 );
buf ( n76111 , n76110 );
buf ( n76112 , n68634 );
not ( n76113 , n69059 );
not ( n76114 , n70139 );
or ( n76115 , n76113 , n76114 );
nand ( n76116 , n70859 , n68661 );
nand ( n76117 , n76115 , n76116 );
buf ( n76118 , n76117 );
buf ( n76119 , 1'b0 );
not ( n76120 , n68838 );
buf ( n9982 , n76120 );
buf ( n9983 , n68634 );
not ( n76123 , n69025 );
not ( n76124 , n70139 );
or ( n76125 , n76123 , n76124 );
nand ( n76126 , n70859 , n2523 );
nand ( n76127 , n76125 , n76126 );
buf ( n76128 , n76127 );
buf ( n76129 , 1'b0 );
not ( n76130 , n68838 );
buf ( n76131 , n76130 );
buf ( n76132 , n68634 );
not ( n76133 , n69083 );
not ( n76134 , n70139 );
or ( n76135 , n76133 , n76134 );
nand ( n76136 , n70859 , n2524 );
nand ( n76137 , n76135 , n76136 );
buf ( n76138 , n76137 );
buf ( n76139 , 1'b0 );
not ( n76140 , n68838 );
buf ( n76141 , n76140 );
buf ( n76142 , n68634 );
not ( n76143 , n69072 );
not ( n76144 , n70139 );
or ( n76145 , n76143 , n76144 );
nand ( n76146 , n70859 , n68664 );
nand ( n76147 , n76145 , n76146 );
buf ( n10009 , n76147 );
buf ( n10010 , 1'b0 );
not ( n76150 , n68838 );
buf ( n76151 , n76150 );
buf ( n76152 , n68634 );
not ( n76153 , n69230 );
or ( n76154 , n71992 , n76153 );
nand ( n76155 , n70859 , n68636 );
nand ( n76156 , n76154 , n76155 );
buf ( n10018 , n76156 );
buf ( n10019 , 1'b0 );
not ( n76159 , n68838 );
buf ( n76160 , n76159 );
buf ( n76161 , n68634 );
not ( n76162 , n69400 );
or ( n76163 , n76162 , n71992 );
nand ( n76164 , n70859 , n2498 );
nand ( n76165 , n76163 , n76164 );
buf ( n76166 , n76165 );
buf ( n76167 , 1'b0 );
not ( n76168 , n68838 );
buf ( n76169 , n76168 );
buf ( n76170 , n68634 );
not ( n76171 , n69095 );
not ( n76172 , n70139 );
or ( n76173 , n76171 , n76172 );
nand ( n76174 , n70859 , n68665 );
nand ( n76175 , n76173 , n76174 );
buf ( n76176 , n76175 );
buf ( n76177 , 1'b0 );
not ( n76178 , n68838 );
buf ( n76179 , n76178 );
buf ( n76180 , n68634 );
not ( n76181 , n69409 );
or ( n76182 , n71992 , n76181 );
nand ( n76183 , n70859 , n2499 );
nand ( n76184 , n76182 , n76183 );
buf ( n76185 , n76184 );
buf ( n76186 , 1'b0 );
not ( n76187 , n68838 );
buf ( n10049 , n76187 );
buf ( n10050 , n68634 );
not ( n76190 , n69352 );
or ( n76191 , n71992 , n76190 );
not ( n76192 , n2500 );
or ( n76193 , n72071 , n76192 );
nand ( n76194 , n76191 , n76193 );
buf ( n76195 , n76194 );
buf ( n76196 , 1'b0 );
not ( n76197 , n68838 );
buf ( n10059 , n76197 );
buf ( n76199 , n68634 );
not ( n76200 , n69338 );
or ( n76201 , n71992 , n76200 );
not ( n76202 , n2501 );
or ( n76203 , n72071 , n76202 );
nand ( n76204 , n76201 , n76203 );
buf ( n10066 , n76204 );
buf ( n10067 , 1'b0 );
not ( n76207 , n68838 );
buf ( n10069 , n76207 );
buf ( n10070 , n68634 );
not ( n76210 , n69324 );
or ( n76211 , n71992 , n76210 );
not ( n76212 , n2502 );
or ( n76213 , n72071 , n76212 );
nand ( n76214 , n76211 , n76213 );
buf ( n76215 , n76214 );
buf ( n76216 , 1'b0 );
not ( n76217 , n68838 );
buf ( n76218 , n76217 );
buf ( n76219 , n68634 );
not ( n76220 , n69298 );
not ( n76221 , n70139 );
or ( n76222 , n76220 , n76221 );
nand ( n76223 , n70859 , n2503 );
nand ( n76224 , n76222 , n76223 );
buf ( n76225 , n76224 );
buf ( n76226 , 1'b0 );
not ( n76227 , n68838 );
buf ( n10089 , n76227 );
buf ( n76229 , n68634 );
not ( n76230 , n69311 );
or ( n76231 , n71992 , n76230 );
not ( n76232 , n2504 );
or ( n76233 , n72071 , n76232 );
nand ( n76234 , n76231 , n76233 );
buf ( n76235 , n76234 );
buf ( n76236 , 1'b0 );
not ( n76237 , n68838 );
buf ( n10099 , n76237 );
buf ( n10100 , n68634 );
not ( n76240 , n69289 );
not ( n76241 , n70139 );
or ( n76242 , n76240 , n76241 );
nand ( n76243 , n70859 , n68644 );
nand ( n76244 , n76242 , n76243 );
buf ( n76245 , n76244 );
buf ( n76246 , 1'b0 );
not ( n76247 , n68838 );
buf ( n76248 , n76247 );
buf ( n76249 , n68634 );
not ( n76250 , n69277 );
or ( n76251 , n71992 , n76250 );
not ( n76252 , n68645 );
or ( n76253 , n72071 , n76252 );
nand ( n76254 , n76251 , n76253 );
buf ( n76255 , n76254 );
buf ( n76256 , 1'b0 );
not ( n76257 , n68838 );
buf ( n10119 , n76257 );
buf ( n10120 , n68634 );
not ( n76260 , n69265 );
or ( n76261 , n71992 , n76260 );
not ( n76262 , n68646 );
or ( n76263 , n72071 , n76262 );
nand ( n76264 , n76261 , n76263 );
buf ( n10126 , n76264 );
buf ( n10127 , 1'b0 );
not ( n76267 , n68838 );
buf ( n10129 , n76267 );
buf ( n10130 , n68634 );
not ( n76270 , n69256 );
or ( n76271 , n71992 , n76270 );
not ( n76272 , n2508 );
or ( n76273 , n72071 , n76272 );
nand ( n76274 , n76271 , n76273 );
buf ( n10136 , n76274 );
buf ( n10137 , 1'b0 );
not ( n76277 , n68838 );
buf ( n76278 , n76277 );
buf ( n10140 , n68634 );
not ( n76280 , n69106 );
not ( n76281 , n70139 );
or ( n76282 , n76280 , n76281 );
nand ( n76283 , n70859 , n68666 );
nand ( n76284 , n76282 , n76283 );
buf ( n76285 , n76284 );
buf ( n76286 , 1'b0 );
not ( n76287 , n68838 );
buf ( n76288 , n76287 );
buf ( n76289 , n68634 );
not ( n76290 , n69240 );
or ( n76291 , n71992 , n76290 );
not ( n76292 , n2509 );
or ( n76293 , n72071 , n76292 );
nand ( n76294 , n76291 , n76293 );
buf ( n10156 , n76294 );
buf ( n76296 , 1'b0 );
not ( n76297 , n68838 );
buf ( n76298 , n76297 );
buf ( n76299 , n68634 );
not ( n76300 , n68649 );
not ( n76301 , n70859 );
or ( n76302 , n76300 , n76301 );
not ( n76303 , n69157 );
or ( n76304 , n71992 , n76303 );
nand ( n76305 , n76302 , n76304 );
buf ( n76306 , n76305 );
buf ( n76307 , 1'b0 );
not ( n76308 , n68838 );
buf ( n76309 , n76308 );
buf ( n76310 , n68634 );
not ( n76311 , n69176 );
or ( n76312 , n71992 , n76311 );
not ( n76313 , n68650 );
or ( n76314 , n72071 , n76313 );
nand ( n76315 , n76312 , n76314 );
buf ( n76316 , n76315 );
buf ( n76317 , 1'b0 );
not ( n76318 , n68838 );
buf ( n76319 , n76318 );
buf ( n76320 , n68634 );
not ( n76321 , n69187 );
not ( n76322 , n70139 );
or ( n76323 , n76321 , n76322 );
nand ( n76324 , n70859 , n68651 );
nand ( n76325 , n76323 , n76324 );
buf ( n76326 , n76325 );
buf ( n76327 , 1'b0 );
not ( n76328 , n68838 );
buf ( n10190 , n76328 );
buf ( n10191 , n68634 );
not ( n76331 , n68934 );
or ( n76332 , n76331 , n71992 );
nand ( n76333 , n70859 , n2513 );
nand ( n76334 , n76332 , n76333 );
buf ( n10196 , n76334 );
buf ( n10197 , 1'b0 );
not ( n76337 , n68838 );
buf ( n76338 , n76337 );
buf ( n76339 , n68634 );
not ( n76340 , n68961 );
or ( n76341 , n71992 , n76340 );
nand ( n76342 , n70859 , n2514 );
nand ( n76343 , n76341 , n76342 );
buf ( n76344 , n76343 );
buf ( n76345 , 1'b0 );
not ( n76346 , n68838 );
buf ( n76347 , n76346 );
buf ( n76348 , n68634 );
not ( n76349 , n68947 );
or ( n76350 , n71992 , n76349 );
nand ( n76351 , n70859 , n2515 );
nand ( n76352 , n76350 , n76351 );
buf ( n76353 , n76352 );
buf ( n76354 , 1'b0 );
not ( n76355 , n68838 );
buf ( n76356 , n76355 );
buf ( n76357 , n68634 );
not ( n76358 , n68908 );
or ( n76359 , n71992 , n76358 );
nand ( n76360 , n70859 , n2516 );
nand ( n76361 , n76359 , n76360 );
buf ( n10223 , n76361 );
buf ( n10224 , 1'b0 );
not ( n76364 , n68838 );
buf ( n76365 , n76364 );
buf ( n76366 , n68634 );
not ( n76367 , n68977 );
or ( n76368 , n71992 , n76367 );
nand ( n76369 , n70859 , n2517 );
nand ( n76370 , n76368 , n76369 );
buf ( n10232 , n76370 );
buf ( n10233 , 1'b0 );
not ( n76373 , n68838 );
buf ( n76374 , n76373 );
buf ( n76375 , n68634 );
not ( n76376 , n69045 );
or ( n76377 , n71992 , n76376 );
nand ( n76378 , n70859 , n2518 );
nand ( n76379 , n76377 , n76378 );
buf ( n76380 , n76379 );
buf ( n76381 , 1'b0 );
not ( n76382 , n68838 );
buf ( n76383 , n76382 );
buf ( n76384 , n68634 );
not ( n76385 , n2728 );
not ( n76386 , n70139 );
or ( n76387 , n76385 , n76386 );
nand ( n76388 , n70859 , n2528 );
nand ( n76389 , n76387 , n76388 );
buf ( n76390 , n76389 );
buf ( n76391 , 1'b0 );
not ( n76392 , n68838 );
buf ( n76393 , n76392 );
buf ( n76394 , n68634 );
not ( n76395 , n69619 );
not ( n76396 , n76395 );
not ( n76397 , n69947 );
nand ( n76398 , n76397 , n73902 );
not ( n76399 , n76398 );
or ( n76400 , n76396 , n76399 );
not ( n76401 , n76398 );
not ( n76402 , n76401 );
and ( n76403 , n69553 , n69543 );
and ( n76404 , n76403 , n69531 , n69519 );
nand ( n76405 , n69470 , n69451 , n69435 , n69471 );
nand ( n76406 , n69487 , n69502 );
nor ( n76407 , n76405 , n76406 );
nand ( n76408 , n76404 , n76407 );
not ( n76409 , n76408 );
and ( n76410 , n69587 , n69576 );
and ( n76411 , n76410 , n69599 );
nand ( n76412 , n76409 , n76411 );
not ( n76413 , n69613 );
xor ( n76414 , n76412 , n76413 );
not ( n76415 , n76414 );
or ( n76416 , n76402 , n76415 );
nand ( n76417 , n76400 , n76416 );
not ( n76418 , n70238 );
nor ( n76419 , n76417 , n76418 );
not ( n76420 , n69599 );
nand ( n76421 , n76404 , n76407 , n76410 );
not ( n76422 , n76421 );
or ( n76423 , n76420 , n76422 );
or ( n76424 , n76421 , n69599 );
nand ( n76425 , n76423 , n76424 );
not ( n76426 , n76425 );
or ( n76427 , n76398 , n76426 );
nand ( n76428 , n76398 , n69981 );
nand ( n76429 , n76427 , n76428 );
not ( n76430 , n70327 );
nor ( n76431 , n76429 , n76430 );
nor ( n76432 , n76419 , n76431 );
not ( n76433 , n70296 );
and ( n76434 , n76403 , n69531 , n69519 );
nand ( n76435 , n76434 , n76407 , n69587 );
xnor ( n76436 , n76435 , n69576 );
not ( n76437 , n76436 );
or ( n76438 , n76398 , n76437 );
nand ( n76439 , n76398 , n70098 );
nand ( n76440 , n76438 , n76439 );
nor ( n76441 , n76433 , n76440 );
not ( n76442 , n70308 );
not ( n76443 , n69990 );
not ( n76444 , n76398 );
not ( n76445 , n76444 );
not ( n76446 , n76445 );
or ( n76447 , n76443 , n76446 );
not ( n76448 , n69587 );
not ( n76449 , n76408 );
or ( n76450 , n76448 , n76449 );
or ( n76451 , n76408 , n69587 );
nand ( n76452 , n76450 , n76451 );
not ( n76453 , n76452 );
or ( n76454 , n76398 , n76453 );
nand ( n76455 , n76447 , n76454 );
nor ( n76456 , n76442 , n76455 );
nor ( n76457 , n76441 , n76456 );
and ( n76458 , n76432 , n76457 );
not ( n76459 , n70378 );
not ( n76460 , n76459 );
not ( n76461 , n70082 );
not ( n76462 , n76398 );
or ( n76463 , n76461 , n76462 );
not ( n76464 , n76401 );
xor ( n76465 , n69553 , n76407 );
not ( n76466 , n76465 );
or ( n76467 , n76464 , n76466 );
nand ( n76468 , n76463 , n76467 );
not ( n76469 , n76468 );
or ( n76470 , n76460 , n76469 );
not ( n76471 , n70263 );
not ( n76472 , n69543 );
nand ( n76473 , n76407 , n69553 );
not ( n76474 , n76473 );
or ( n76475 , n76472 , n76474 );
or ( n76476 , n76473 , n69543 );
nand ( n76477 , n76475 , n76476 );
not ( n76478 , n76477 );
or ( n76479 , n76398 , n76478 );
nand ( n76480 , n76398 , n70007 );
nand ( n76481 , n76479 , n76480 );
nand ( n76482 , n76471 , n76481 );
nand ( n76483 , n76470 , n76482 );
not ( n76484 , n76481 );
nand ( n76485 , n76484 , n70263 );
nand ( n76486 , n76483 , n76485 );
not ( n76487 , n70253 );
not ( n76488 , n70013 );
not ( n76489 , n76398 );
or ( n76490 , n76488 , n76489 );
not ( n76491 , n69531 );
nand ( n76492 , n76407 , n76403 );
not ( n76493 , n76492 );
or ( n76494 , n76491 , n76493 );
or ( n76495 , n76492 , n69531 );
nand ( n76496 , n76494 , n76495 );
not ( n76497 , n76496 );
or ( n76498 , n76402 , n76497 );
nand ( n76499 , n76490 , n76498 );
not ( n76500 , n76499 );
not ( n76501 , n76500 );
or ( n76502 , n76487 , n76501 );
not ( n76503 , n69519 );
nand ( n76504 , n76407 , n76403 , n69531 );
not ( n76505 , n76504 );
or ( n76506 , n76503 , n76505 );
or ( n76507 , n76504 , n69519 );
nand ( n76508 , n76506 , n76507 );
not ( n76509 , n76508 );
or ( n76510 , n76398 , n76509 );
not ( n76511 , n76398 );
not ( n76512 , n76511 );
not ( n76513 , n71529 );
nand ( n76514 , n76512 , n76513 );
nand ( n76515 , n76510 , n76514 );
not ( n76516 , n70273 );
nor ( n76517 , n76515 , n76516 );
not ( n76518 , n76517 );
nand ( n76519 , n76502 , n76518 );
or ( n76520 , n76486 , n76519 );
not ( n76521 , n70253 );
nand ( n76522 , n76521 , n76499 );
or ( n76523 , n76517 , n76522 );
not ( n76524 , n76515 );
or ( n76525 , n76524 , n70273 );
nand ( n76526 , n76523 , n76525 );
not ( n76527 , n76526 );
nand ( n76528 , n76520 , n76527 );
and ( n76529 , n76458 , n76528 );
not ( n76530 , n76432 );
not ( n76531 , n70308 );
nand ( n76532 , n76531 , n76455 );
or ( n76533 , n76441 , n76532 );
not ( n76534 , n76440 );
or ( n76535 , n76534 , n70296 );
nand ( n76536 , n76533 , n76535 );
not ( n76537 , n76536 );
or ( n76538 , n76530 , n76537 );
not ( n76539 , n76419 );
nand ( n76540 , n76429 , n76430 );
not ( n76541 , n76540 );
and ( n76542 , n76539 , n76541 );
and ( n76543 , n76417 , n76418 );
nor ( n76544 , n76542 , n76543 );
nand ( n76545 , n76538 , n76544 );
nor ( n76546 , n76529 , n76545 );
not ( n76547 , n70378 );
not ( n76548 , n76468 );
not ( n76549 , n76548 );
or ( n76550 , n76547 , n76549 );
nand ( n76551 , n76550 , n76485 );
nor ( n76552 , n76551 , n76519 );
not ( n76553 , n70024 );
not ( n76554 , n76398 );
or ( n76555 , n76553 , n76554 );
not ( n76556 , n76398 );
not ( n76557 , n69502 );
nand ( n76558 , n69451 , n69471 );
not ( n76559 , n76558 );
nand ( n76560 , n76559 , n69487 );
not ( n76561 , n76560 );
or ( n76562 , n76557 , n76561 );
or ( n76563 , n76560 , n69502 );
nand ( n76564 , n76562 , n76563 );
nand ( n76565 , n76556 , n76564 );
nand ( n76566 , n76555 , n76565 );
not ( n76567 , n70432 );
nor ( n76568 , n76566 , n76567 );
not ( n76569 , n72302 );
not ( n76570 , n69487 );
not ( n76571 , n76558 );
or ( n76572 , n76570 , n76571 );
or ( n76573 , n76558 , n69487 );
nand ( n76574 , n76572 , n76573 );
not ( n76575 , n76574 );
or ( n76576 , n76398 , n76575 );
nand ( n76577 , n76512 , n70038 );
nand ( n76578 , n76576 , n76577 );
nor ( n76579 , n76569 , n76578 );
nor ( n76580 , n76568 , n76579 );
not ( n76581 , n69470 );
not ( n76582 , n76406 );
nand ( n76583 , n76582 , n76559 , n69435 );
not ( n76584 , n76583 );
or ( n76585 , n76581 , n76584 );
or ( n76586 , n76583 , n69470 );
nand ( n76587 , n76585 , n76586 );
not ( n76588 , n76587 );
or ( n76589 , n76398 , n76588 );
nand ( n76590 , n76512 , n70090 );
nand ( n76591 , n76589 , n76590 );
not ( n76592 , n70388 );
nor ( n76593 , n76591 , n76592 );
not ( n76594 , n70031 );
not ( n76595 , n76398 );
or ( n76596 , n76594 , n76595 );
not ( n76597 , n76444 );
not ( n76598 , n69435 );
or ( n76599 , n76558 , n76406 );
not ( n76600 , n76599 );
or ( n76601 , n76598 , n76600 );
or ( n76602 , n76599 , n69435 );
nand ( n76603 , n76601 , n76602 );
not ( n76604 , n76603 );
or ( n76605 , n76597 , n76604 );
nand ( n76606 , n76596 , n76605 );
not ( n76607 , n70477 );
nor ( n76608 , n76606 , n76607 );
nor ( n76609 , n76593 , n76608 );
not ( n76610 , n70420 );
not ( n76611 , n76610 );
not ( n76612 , n69451 );
not ( n76613 , n69471 );
and ( n76614 , n76612 , n76613 );
nor ( n76615 , n76614 , n76559 );
not ( n76616 , n76615 );
or ( n76617 , n76398 , n76616 );
nand ( n76618 , n76512 , n70040 );
nand ( n76619 , n76617 , n76618 );
not ( n76620 , n76619 );
or ( n76621 , n76611 , n76620 );
or ( n76622 , n76619 , n76610 );
not ( n76623 , n70053 );
nand ( n76624 , n76623 , n70503 );
not ( n76625 , n69967 );
nand ( n76626 , n76625 , n70522 );
and ( n76627 , n76624 , n76626 );
not ( n76628 , n70503 );
and ( n76629 , n70053 , n76628 );
nor ( n76630 , n76627 , n76629 );
not ( n76631 , n70073 );
and ( n76632 , n76631 , n70459 );
or ( n76633 , n76630 , n76632 );
or ( n76634 , n76631 , n70459 );
nand ( n76635 , n76633 , n76634 );
nand ( n76636 , n76622 , n76635 );
nand ( n76637 , n76621 , n76636 );
nand ( n76638 , n76580 , n76609 , n76637 );
not ( n76639 , n72302 );
nand ( n76640 , n76639 , n76578 );
not ( n76641 , n70432 );
nand ( n76642 , n76641 , n76566 );
and ( n76643 , n76640 , n76642 );
nor ( n76644 , n76643 , n76568 );
nand ( n76645 , n76644 , n76609 );
nand ( n76646 , n76606 , n76607 );
nor ( n76647 , n76593 , n76646 );
and ( n76648 , n76591 , n76592 );
nor ( n76649 , n76647 , n76648 );
nand ( n76650 , n76638 , n76645 , n76649 );
nand ( n76651 , n76552 , n76458 , n76650 );
nand ( n76652 , n76546 , n76651 );
and ( n76653 , n69599 , n69613 );
nand ( n76654 , n76410 , n76653 );
nor ( n76655 , n76408 , n76654 );
nand ( n76656 , n69655 , n69641 );
nand ( n76657 , n69896 , n69769 );
nor ( n76658 , n76656 , n76657 );
and ( n76659 , n69822 , n69871 , n69804 , n69792 );
nand ( n76660 , n76658 , n76659 );
nand ( n76661 , n69932 , n69850 );
nand ( n76662 , n69685 , n69706 );
nor ( n76663 , n76661 , n76662 );
not ( n76664 , n72628 );
nand ( n76665 , n76663 , n76664 );
nor ( n76666 , n76660 , n76665 );
nand ( n76667 , n76655 , n76666 );
not ( n76668 , n69743 );
and ( n76669 , n76667 , n76668 );
not ( n76670 , n76667 );
and ( n76671 , n76670 , n69743 );
nor ( n76672 , n76669 , n76671 );
not ( n76673 , n76672 );
or ( n76674 , n76445 , n76673 );
nand ( n76675 , n76398 , n72463 );
nand ( n76676 , n76674 , n76675 );
not ( n76677 , n76676 );
nand ( n76678 , n76677 , n73916 );
not ( n76679 , n76663 );
nand ( n76680 , n76658 , n76659 );
nor ( n76681 , n76679 , n76680 );
nand ( n76682 , n76655 , n76681 );
not ( n76683 , n76664 );
and ( n76684 , n76682 , n76683 );
not ( n76685 , n76682 );
and ( n76686 , n76685 , n76664 );
nor ( n76687 , n76684 , n76686 );
not ( n76688 , n76687 );
or ( n76689 , n76398 , n76688 );
nand ( n76690 , n76512 , n72452 );
nand ( n76691 , n76689 , n76690 );
not ( n76692 , n76691 );
nand ( n76693 , n76692 , n72626 );
nand ( n76694 , n76678 , n76693 );
not ( n76695 , n73914 );
nand ( n76696 , n76664 , n69743 );
not ( n76697 , n76696 );
nand ( n76698 , n76697 , n76663 );
nor ( n76699 , n76680 , n76698 );
nand ( n76700 , n76655 , n76699 );
and ( n76701 , n76700 , n69908 );
not ( n76702 , n76700 );
not ( n76703 , n69908 );
and ( n76704 , n76702 , n76703 );
nor ( n76705 , n76701 , n76704 );
not ( n76706 , n76705 );
or ( n76707 , n76398 , n76706 );
nand ( n76708 , n76398 , n73902 );
nand ( n76709 , n76707 , n76708 );
not ( n76710 , n76709 );
not ( n76711 , n76710 );
or ( n76712 , n76695 , n76711 );
nor ( n76713 , n76696 , n69908 );
nand ( n76714 , n76663 , n76713 );
nor ( n76715 , n76680 , n76714 );
nand ( n76716 , n76655 , n76715 );
not ( n76717 , n69942 );
and ( n76718 , n76717 , n76703 );
not ( n76719 , n76717 );
and ( n76720 , n76719 , n69908 );
nor ( n76721 , n76718 , n76720 );
xor ( n76722 , n76716 , n76721 );
not ( n76723 , n76722 );
not ( n76724 , n76398 );
not ( n76725 , n76724 );
or ( n76726 , n76723 , n76725 );
not ( n76727 , n69947 );
nand ( n76728 , n76726 , n76727 );
not ( n76729 , n73912 );
nand ( n76730 , n76728 , n76729 );
nand ( n76731 , n76712 , n76730 );
nor ( n76732 , n76694 , n76731 );
not ( n76733 , n76661 );
nand ( n76734 , n76733 , n69685 );
nor ( n76735 , n76660 , n76734 );
nand ( n76736 , n76655 , n76735 );
not ( n76737 , n69706 );
and ( n76738 , n76736 , n76737 );
not ( n76739 , n76736 );
and ( n76740 , n76739 , n69706 );
nor ( n76741 , n76738 , n76740 );
not ( n76742 , n76741 );
or ( n76743 , n76597 , n76742 );
nand ( n76744 , n76398 , n71763 );
nand ( n76745 , n76743 , n76744 );
not ( n76746 , n72815 );
nor ( n76747 , n76745 , n76746 );
not ( n76748 , n71779 );
not ( n76749 , n76748 );
not ( n76750 , n76512 );
or ( n76751 , n76749 , n76750 );
nor ( n76752 , n76660 , n76661 );
nand ( n76753 , n76655 , n76752 );
not ( n76754 , n69685 );
and ( n76755 , n76753 , n76754 );
not ( n76756 , n76753 );
and ( n76757 , n76756 , n69685 );
nor ( n76758 , n76755 , n76757 );
not ( n76759 , n76758 );
or ( n76760 , n76597 , n76759 );
nand ( n76761 , n76751 , n76760 );
not ( n76762 , n72534 );
nor ( n76763 , n76761 , n76762 );
nor ( n76764 , n76747 , n76763 );
not ( n76765 , n76764 );
not ( n76766 , n72557 );
not ( n76767 , n76680 );
nand ( n76768 , n76767 , n76655 );
not ( n76769 , n69932 );
and ( n76770 , n76768 , n76769 );
not ( n76771 , n76768 );
and ( n76772 , n76771 , n69932 );
nor ( n76773 , n76770 , n76772 );
not ( n76774 , n76773 );
or ( n76775 , n76398 , n76774 );
nand ( n76776 , n76398 , n71814 );
nand ( n76777 , n76775 , n76776 );
not ( n76778 , n76777 );
not ( n76779 , n76778 );
or ( n76780 , n76766 , n76779 );
not ( n76781 , n71798 );
not ( n76782 , n76781 );
not ( n76783 , n76398 );
or ( n76784 , n76782 , n76783 );
nor ( n76785 , n76660 , n76769 );
nand ( n76786 , n76655 , n76785 );
not ( n76787 , n69850 );
and ( n76788 , n76786 , n76787 );
not ( n76789 , n76786 );
and ( n76790 , n76789 , n69850 );
nor ( n76791 , n76788 , n76790 );
not ( n76792 , n76791 );
or ( n76793 , n76398 , n76792 );
nand ( n76794 , n76784 , n76793 );
not ( n76795 , n72544 );
nor ( n76796 , n76794 , n76795 );
not ( n76797 , n76796 );
nand ( n76798 , n76780 , n76797 );
nor ( n76799 , n76765 , n76798 );
nand ( n76800 , n76732 , n76799 );
nand ( n76801 , n69804 , n69822 );
nor ( n76802 , n76656 , n76801 );
nand ( n76803 , n69896 , n69871 );
not ( n76804 , n69792 );
nor ( n76805 , n76803 , n76804 );
and ( n76806 , n76802 , n76805 );
nand ( n76807 , n76655 , n76806 );
not ( n76808 , n69769 );
and ( n76809 , n76807 , n76808 );
not ( n76810 , n76807 );
and ( n76811 , n76810 , n69769 );
nor ( n76812 , n76809 , n76811 );
not ( n76813 , n76812 );
or ( n76814 , n76597 , n76813 );
not ( n76815 , n71833 );
nand ( n76816 , n76398 , n76815 );
nand ( n76817 , n76814 , n76816 );
not ( n76818 , n72510 );
nor ( n76819 , n76817 , n76818 );
not ( n76820 , n72499 );
not ( n76821 , n71852 );
not ( n76822 , n76445 );
or ( n76823 , n76821 , n76822 );
not ( n76824 , n76803 );
and ( n76825 , n76802 , n76824 );
nand ( n76826 , n76655 , n76825 );
and ( n76827 , n76826 , n76804 );
not ( n76828 , n76826 );
and ( n76829 , n76828 , n69792 );
nor ( n76830 , n76827 , n76829 );
not ( n76831 , n76830 );
or ( n76832 , n76398 , n76831 );
nand ( n76833 , n76823 , n76832 );
nor ( n76834 , n76820 , n76833 );
nor ( n76835 , n76819 , n76834 );
not ( n76836 , n71869 );
not ( n76837 , n76398 );
or ( n76838 , n76836 , n76837 );
and ( n76839 , n76802 , n69871 );
nand ( n76840 , n76655 , n76839 );
not ( n76841 , n69896 );
and ( n76842 , n76840 , n76841 );
not ( n76843 , n76840 );
and ( n76844 , n76843 , n69896 );
nor ( n76845 , n76842 , n76844 );
not ( n76846 , n76845 );
or ( n76847 , n76464 , n76846 );
nand ( n76848 , n76838 , n76847 );
not ( n76849 , n72475 );
nor ( n76850 , n76848 , n76849 );
not ( n76851 , n71037 );
not ( n76852 , n76398 );
or ( n76853 , n76851 , n76852 );
nand ( n76854 , n76655 , n76802 );
not ( n76855 , n69871 );
and ( n76856 , n76854 , n76855 );
not ( n76857 , n76854 );
and ( n76858 , n76857 , n69871 );
nor ( n76859 , n76856 , n76858 );
not ( n76860 , n76859 );
or ( n76861 , n76402 , n76860 );
nand ( n76862 , n76853 , n76861 );
not ( n76863 , n72485 );
nor ( n76864 , n76862 , n76863 );
nor ( n76865 , n76850 , n76864 );
and ( n76866 , n76835 , n76865 );
not ( n76867 , n70225 );
not ( n76868 , n69977 );
not ( n76869 , n76398 );
or ( n76870 , n76868 , n76869 );
xor ( n76871 , n69641 , n76655 );
not ( n76872 , n76871 );
or ( n76873 , n76398 , n76872 );
nand ( n76874 , n76870 , n76873 );
not ( n76875 , n76874 );
not ( n76876 , n76875 );
or ( n76877 , n76867 , n76876 );
nand ( n76878 , n76655 , n69641 );
not ( n76879 , n69655 );
and ( n76880 , n76878 , n76879 );
not ( n76881 , n76878 );
and ( n76882 , n76881 , n69655 );
nor ( n76883 , n76880 , n76882 );
not ( n76884 , n76883 );
or ( n76885 , n76398 , n76884 );
nand ( n76886 , n76445 , n69660 );
nand ( n76887 , n76885 , n76886 );
not ( n76888 , n76887 );
nand ( n76889 , n76888 , n71074 );
nand ( n76890 , n76877 , n76889 );
not ( n76891 , n71092 );
not ( n76892 , n71047 );
not ( n76893 , n76398 );
or ( n76894 , n76892 , n76893 );
not ( n76895 , n76656 );
nand ( n76896 , n76895 , n76655 );
not ( n76897 , n69822 );
and ( n76898 , n76896 , n76897 );
not ( n76899 , n76896 );
and ( n76900 , n76899 , n69822 );
nor ( n76901 , n76898 , n76900 );
not ( n76902 , n76901 );
or ( n76903 , n76402 , n76902 );
nand ( n76904 , n76894 , n76903 );
not ( n76905 , n76904 );
not ( n76906 , n76905 );
or ( n76907 , n76891 , n76906 );
nor ( n76908 , n76656 , n76897 );
nand ( n76909 , n76655 , n76908 );
xnor ( n76910 , n76909 , n69804 );
not ( n76911 , n76910 );
not ( n76912 , n76401 );
or ( n76913 , n76911 , n76912 );
not ( n76914 , n76398 );
not ( n76915 , n71058 );
or ( n76916 , n76914 , n76915 );
nand ( n76917 , n76913 , n76916 );
not ( n76918 , n71122 );
nor ( n76919 , n76917 , n76918 );
not ( n76920 , n76919 );
nand ( n76921 , n76907 , n76920 );
nor ( n76922 , n76890 , n76921 );
nand ( n76923 , n76866 , n76922 );
nor ( n76924 , n76800 , n76923 );
and ( n76925 , n76652 , n76924 );
not ( n76926 , n71074 );
nand ( n76927 , n76926 , n76887 );
not ( n76928 , n76927 );
not ( n76929 , n70225 );
nand ( n76930 , n76929 , n76874 );
not ( n76931 , n76930 );
or ( n76932 , n76928 , n76931 );
nand ( n76933 , n76932 , n76889 );
or ( n76934 , n76921 , n76933 );
not ( n76935 , n71092 );
nand ( n76936 , n76935 , n76904 );
or ( n76937 , n76919 , n76936 );
nand ( n76938 , n76917 , n76918 );
nand ( n76939 , n76937 , n76938 );
not ( n76940 , n76939 );
nand ( n76941 , n76934 , n76940 );
and ( n76942 , n76866 , n76941 );
not ( n76943 , n76835 );
nand ( n76944 , n76862 , n76863 );
or ( n76945 , n76850 , n76944 );
nand ( n76946 , n76848 , n76849 );
nand ( n76947 , n76945 , n76946 );
not ( n76948 , n76947 );
or ( n76949 , n76943 , n76948 );
not ( n76950 , n76819 );
not ( n76951 , n72499 );
nand ( n76952 , n76951 , n76833 );
not ( n76953 , n76952 );
and ( n76954 , n76950 , n76953 );
and ( n76955 , n76817 , n76818 );
nor ( n76956 , n76954 , n76955 );
nand ( n76957 , n76949 , n76956 );
nor ( n76958 , n76942 , n76957 );
or ( n76959 , n76958 , n76800 );
not ( n76960 , n76764 );
not ( n76961 , n72557 );
nand ( n76962 , n76961 , n76777 );
or ( n76963 , n76796 , n76962 );
nand ( n76964 , n76794 , n76795 );
nand ( n76965 , n76963 , n76964 );
not ( n76966 , n76965 );
or ( n76967 , n76960 , n76966 );
not ( n76968 , n76747 );
nand ( n76969 , n76761 , n76762 );
not ( n76970 , n76969 );
and ( n76971 , n76968 , n76970 );
and ( n76972 , n76745 , n76746 );
nor ( n76973 , n76971 , n76972 );
nand ( n76974 , n76967 , n76973 );
and ( n76975 , n76974 , n76732 );
not ( n76976 , n76691 );
nor ( n76977 , n76976 , n72626 );
and ( n76978 , n76678 , n76977 );
not ( n76979 , n76676 );
nor ( n76980 , n76979 , n73916 );
nor ( n76981 , n76978 , n76980 );
or ( n76982 , n76981 , n76731 );
nor ( n76983 , n76710 , n73914 );
and ( n76984 , n76983 , n76730 );
nor ( n76985 , n76728 , n76729 );
nor ( n76986 , n76984 , n76985 );
nand ( n76987 , n76982 , n76986 );
nor ( n76988 , n76975 , n76987 );
nand ( n76989 , n76959 , n76988 );
nor ( n76990 , n76925 , n76989 );
not ( n76991 , n76990 );
not ( n76992 , n72499 );
not ( n76993 , n76992 );
not ( n76994 , n71852 );
or ( n76995 , n76993 , n76994 );
not ( n76996 , n72510 );
nand ( n76997 , n76815 , n76996 );
nand ( n76998 , n76995 , n76997 );
not ( n76999 , n72485 );
not ( n77000 , n76999 );
not ( n77001 , n71037 );
or ( n77002 , n77000 , n77001 );
not ( n77003 , n72475 );
nand ( n77004 , n71869 , n77003 );
nand ( n77005 , n77002 , n77004 );
nor ( n77006 , n76998 , n77005 );
not ( n77007 , n71092 );
not ( n77008 , n77007 );
not ( n77009 , n71047 );
or ( n77010 , n77008 , n77009 );
not ( n77011 , n71122 );
nand ( n77012 , n71058 , n77011 );
nand ( n77013 , n77010 , n77012 );
not ( n77014 , n71074 );
not ( n77015 , n69660 );
not ( n77016 , n77015 );
or ( n77017 , n77014 , n77016 );
not ( n77018 , n69977 );
nand ( n77019 , n77018 , n70225 );
nand ( n77020 , n77017 , n77019 );
not ( n77021 , n71074 );
nand ( n77022 , n77021 , n69660 );
nand ( n77023 , n77020 , n77022 );
or ( n77024 , n77013 , n77023 );
nor ( n77025 , n71047 , n77007 );
and ( n77026 , n77012 , n77025 );
nor ( n77027 , n71058 , n77011 );
nor ( n77028 , n77026 , n77027 );
nand ( n77029 , n77024 , n77028 );
and ( n77030 , n77006 , n77029 );
nor ( n77031 , n71037 , n76999 );
and ( n77032 , n77004 , n77031 );
nor ( n77033 , n71869 , n77003 );
nor ( n77034 , n77032 , n77033 );
or ( n77035 , n77034 , n76998 );
nor ( n77036 , n71852 , n76992 );
and ( n77037 , n76997 , n77036 );
nor ( n77038 , n76815 , n76996 );
nor ( n77039 , n77037 , n77038 );
nand ( n77040 , n77035 , n77039 );
nor ( n77041 , n77030 , n77040 );
not ( n77042 , n72626 );
not ( n77043 , n77042 );
not ( n77044 , n72452 );
or ( n77045 , n77043 , n77044 );
not ( n77046 , n73916 );
nand ( n77047 , n77046 , n72463 );
nand ( n77048 , n77045 , n77047 );
not ( n77049 , n73914 );
not ( n77050 , n77049 );
not ( n77051 , n73902 );
or ( n77052 , n77050 , n77051 );
not ( n77053 , n69947 );
nand ( n77054 , n77053 , n73912 );
nand ( n77055 , n77052 , n77054 );
nor ( n77056 , n77048 , n77055 );
not ( n77057 , n72534 );
not ( n77058 , n77057 );
not ( n77059 , n76748 );
or ( n77060 , n77058 , n77059 );
not ( n77061 , n72815 );
nand ( n77062 , n71763 , n77061 );
nand ( n77063 , n77060 , n77062 );
not ( n77064 , n72557 );
not ( n77065 , n77064 );
not ( n77066 , n71814 );
or ( n77067 , n77065 , n77066 );
not ( n77068 , n72544 );
nand ( n77069 , n76781 , n77068 );
nand ( n77070 , n77067 , n77069 );
nor ( n77071 , n77063 , n77070 );
nand ( n77072 , n77056 , n77071 );
or ( n77073 , n77041 , n77072 );
nor ( n77074 , n76781 , n77068 );
nor ( n77075 , n71814 , n77064 );
or ( n77076 , n77074 , n77075 );
nand ( n77077 , n77076 , n77069 );
or ( n77078 , n77063 , n77077 );
nor ( n77079 , n76748 , n77057 );
and ( n77080 , n77062 , n77079 );
nor ( n77081 , n71763 , n77061 );
nor ( n77082 , n77080 , n77081 );
nand ( n77083 , n77078 , n77082 );
and ( n77084 , n77056 , n77083 );
not ( n77085 , n72463 );
not ( n77086 , n73916 );
not ( n77087 , n77086 );
and ( n77088 , n77085 , n77087 );
nor ( n77089 , n72452 , n77042 );
and ( n77090 , n77047 , n77089 );
nor ( n77091 , n77088 , n77090 );
or ( n77092 , n77091 , n77055 );
nor ( n77093 , n73902 , n77049 );
and ( n77094 , n77054 , n77093 );
not ( n77095 , n69947 );
nor ( n77096 , n77095 , n73912 );
nor ( n77097 , n77094 , n77096 );
nand ( n77098 , n77092 , n77097 );
nor ( n77099 , n77084 , n77098 );
nand ( n77100 , n77073 , n77099 );
not ( n77101 , n70225 );
not ( n77102 , n77101 );
not ( n77103 , n69977 );
or ( n77104 , n77102 , n77103 );
nand ( n77105 , n77104 , n77022 );
nor ( n77106 , n77013 , n77105 );
nand ( n77107 , n77006 , n77106 );
not ( n77108 , n70327 );
not ( n77109 , n77108 );
not ( n77110 , n69981 );
or ( n77111 , n77109 , n77110 );
not ( n77112 , n70238 );
nand ( n77113 , n77112 , n76395 );
nand ( n77114 , n77111 , n77113 );
not ( n77115 , n70308 );
not ( n77116 , n77115 );
not ( n77117 , n69990 );
or ( n77118 , n77116 , n77117 );
not ( n77119 , n70296 );
nand ( n77120 , n77119 , n70098 );
nand ( n77121 , n77118 , n77120 );
nor ( n77122 , n77114 , n77121 );
not ( n77123 , n70253 );
not ( n77124 , n77123 );
not ( n77125 , n70013 );
or ( n77126 , n77124 , n77125 );
not ( n77127 , n71529 );
not ( n77128 , n70273 );
nand ( n77129 , n77127 , n77128 );
nand ( n77130 , n77126 , n77129 );
not ( n77131 , n70378 );
not ( n77132 , n77131 );
not ( n77133 , n70082 );
or ( n77134 , n77132 , n77133 );
not ( n77135 , n70263 );
nand ( n77136 , n77135 , n70007 );
nand ( n77137 , n77134 , n77136 );
nor ( n77138 , n77130 , n77137 );
not ( n77139 , n70388 );
nand ( n77140 , n70090 , n77139 );
not ( n77141 , n70477 );
nand ( n77142 , n77141 , n70031 );
and ( n77143 , n77140 , n77142 );
not ( n77144 , n70432 );
nand ( n77145 , n77144 , n70024 );
not ( n77146 , n70817 );
not ( n77147 , n77146 );
nand ( n77148 , n77147 , n70038 );
and ( n77149 , n77145 , n77148 );
not ( n77150 , n70420 );
nand ( n77151 , n77150 , n70040 );
not ( n77152 , n69967 );
nor ( n77153 , n77152 , n70522 );
not ( n77154 , n70053 );
nor ( n77155 , n77154 , n70503 );
or ( n77156 , n77153 , n77155 );
not ( n77157 , n70503 );
or ( n77158 , n70053 , n77157 );
nand ( n77159 , n77156 , n77158 );
not ( n77160 , n70459 );
nand ( n77161 , n77160 , n70073 );
nand ( n77162 , n77151 , n77159 , n77161 );
not ( n77163 , n70459 );
nor ( n77164 , n77163 , n70073 );
nand ( n77165 , n77151 , n77164 );
not ( n77166 , n70040 );
nand ( n77167 , n77166 , n70420 );
nand ( n77168 , n77162 , n77165 , n77167 );
nand ( n77169 , n77143 , n77149 , n77168 );
not ( n77170 , n77146 );
nor ( n77171 , n77170 , n70038 );
not ( n77172 , n77171 );
not ( n77173 , n77145 );
or ( n77174 , n77172 , n77173 );
not ( n77175 , n70024 );
nand ( n77176 , n77175 , n70432 );
nand ( n77177 , n77174 , n77176 );
nand ( n77178 , n77143 , n77177 );
not ( n77179 , n70477 );
nor ( n77180 , n77179 , n70031 );
and ( n77181 , n77140 , n77180 );
nor ( n77182 , n70090 , n77139 );
nor ( n77183 , n77181 , n77182 );
nand ( n77184 , n77169 , n77178 , n77183 );
and ( n77185 , n77122 , n77138 , n77184 );
not ( n77186 , n77122 );
nor ( n77187 , n70082 , n77131 );
and ( n77188 , n77136 , n77187 );
not ( n77189 , n70007 );
and ( n77190 , n77189 , n70263 );
nor ( n77191 , n77188 , n77190 );
or ( n77192 , n77191 , n77130 );
nor ( n77193 , n70013 , n77123 );
and ( n77194 , n77129 , n77193 );
nor ( n77195 , n77127 , n77128 );
nor ( n77196 , n77194 , n77195 );
nand ( n77197 , n77192 , n77196 );
not ( n77198 , n77197 );
or ( n77199 , n77186 , n77198 );
not ( n77200 , n77114 );
nor ( n77201 , n69990 , n77115 );
not ( n77202 , n77201 );
not ( n77203 , n77120 );
or ( n77204 , n77202 , n77203 );
not ( n77205 , n70098 );
nand ( n77206 , n77205 , n70296 );
nand ( n77207 , n77204 , n77206 );
and ( n77208 , n77200 , n77207 );
nor ( n77209 , n69981 , n77108 );
not ( n77210 , n77209 );
not ( n77211 , n77113 );
or ( n77212 , n77210 , n77211 );
not ( n77213 , n76395 );
nand ( n77214 , n77213 , n70238 );
nand ( n77215 , n77212 , n77214 );
nor ( n77216 , n77208 , n77215 );
nand ( n77217 , n77199 , n77216 );
nor ( n77218 , n77185 , n77217 );
nor ( n77219 , n77107 , n77218 , n77072 );
nor ( n77220 , n77100 , n77219 );
nand ( n77221 , n70196 , n70147 );
or ( n77222 , n77220 , n77221 );
or ( n77223 , n77221 , n70152 );
nand ( n77224 , n77222 , n77223 );
nand ( n77225 , n77224 , n71983 );
not ( n77226 , n70194 );
nor ( n77227 , n77226 , n70188 );
nand ( n77228 , n77227 , n70147 );
nand ( n77229 , n77221 , n77228 );
not ( n77230 , n77229 );
not ( n77231 , n77220 );
or ( n77232 , n77230 , n77231 );
nand ( n77233 , n77232 , n77223 );
nand ( n77234 , n77233 , n70874 );
not ( n77235 , n77220 );
not ( n77236 , n77228 );
nand ( n77237 , n77236 , n71983 );
not ( n77238 , n77237 );
and ( n77239 , n77235 , n77238 );
and ( n77240 , n70202 , n70206 , n70139 );
not ( n77241 , n77240 );
not ( n77242 , n70225 );
nand ( n77243 , n77242 , n69641 );
not ( n77244 , n69641 );
nand ( n77245 , n77244 , n70225 );
nand ( n77246 , n77243 , n77245 );
not ( n77247 , n70238 );
nand ( n77248 , n77247 , n69613 );
and ( n77249 , n77246 , n77248 );
not ( n77250 , n77246 );
not ( n77251 , n77248 );
and ( n77252 , n77250 , n77251 );
nor ( n77253 , n77249 , n77252 );
not ( n77254 , n72557 );
nand ( n77255 , n77254 , n69932 );
not ( n77256 , n69932 );
nand ( n77257 , n77256 , n72557 );
nand ( n77258 , n77255 , n77257 );
not ( n77259 , n72510 );
nand ( n77260 , n77259 , n69769 );
xor ( n77261 , n77258 , n77260 );
nand ( n77262 , n77253 , n77261 );
not ( n77263 , n72626 );
nand ( n77264 , n77263 , n69729 );
not ( n77265 , n69729 );
nand ( n77266 , n77265 , n72626 );
nand ( n77267 , n77264 , n77266 );
not ( n77268 , n72814 );
not ( n77269 , n77268 );
nand ( n77270 , n77269 , n69706 );
xor ( n77271 , n77267 , n77270 );
not ( n77272 , n73916 );
nand ( n77273 , n77272 , n69743 );
not ( n77274 , n77273 );
not ( n77275 , n77274 );
not ( n77276 , n73914 );
nand ( n77277 , n77276 , n69908 );
not ( n77278 , n69908 );
nand ( n77279 , n77278 , n73914 );
nand ( n77280 , n77277 , n77279 );
not ( n77281 , n77280 );
or ( n77282 , n77275 , n77281 );
or ( n77283 , n77280 , n77274 );
nand ( n77284 , n77282 , n77283 );
not ( n77285 , n77277 );
not ( n77286 , n77285 );
xor ( n77287 , n69942 , n73912 );
not ( n77288 , n77287 );
or ( n77289 , n77286 , n77288 );
or ( n77290 , n77287 , n77285 );
nand ( n77291 , n77289 , n77290 );
nand ( n77292 , n77271 , n77284 , n77291 );
nor ( n77293 , n77262 , n77292 );
not ( n77294 , n71122 );
not ( n77295 , n69804 );
not ( n77296 , n77295 );
or ( n77297 , n77294 , n77296 );
not ( n77298 , n71122 );
nand ( n77299 , n77298 , n69804 );
nand ( n77300 , n77297 , n77299 );
not ( n77301 , n77300 );
not ( n77302 , n71092 );
nand ( n77303 , n77302 , n69822 );
not ( n77304 , n77303 );
and ( n77305 , n77301 , n77304 );
and ( n77306 , n77300 , n77303 );
nor ( n77307 , n77305 , n77306 );
not ( n77308 , n71092 );
not ( n77309 , n69822 );
not ( n77310 , n77309 );
or ( n77311 , n77308 , n77310 );
nand ( n77312 , n77311 , n77303 );
not ( n77313 , n71074 );
nand ( n77314 , n77313 , n69655 );
and ( n77315 , n77312 , n77314 );
not ( n77316 , n77312 );
not ( n77317 , n77314 );
and ( n77318 , n77316 , n77317 );
nor ( n77319 , n77315 , n77318 );
not ( n77320 , n69576 );
not ( n77321 , n77320 );
not ( n77322 , n70296 );
or ( n77323 , n77321 , n77322 );
not ( n77324 , n70296 );
nand ( n77325 , n77324 , n69576 );
nand ( n77326 , n77323 , n77325 );
not ( n77327 , n70308 );
nand ( n77328 , n77327 , n69587 );
xor ( n77329 , n77326 , n77328 );
not ( n77330 , n72499 );
nand ( n77331 , n77330 , n69792 );
not ( n77332 , n69792 );
nand ( n77333 , n77332 , n72499 );
nand ( n77334 , n77331 , n77333 );
not ( n77335 , n72475 );
nand ( n77336 , n77335 , n69896 );
xor ( n77337 , n77334 , n77336 );
nand ( n77338 , n77307 , n77319 , n77329 , n77337 );
not ( n77339 , n72544 );
nand ( n77340 , n77339 , n69850 );
not ( n77341 , n69850 );
nand ( n77342 , n77341 , n72544 );
nand ( n77343 , n77340 , n77342 );
xor ( n77344 , n77343 , n77255 );
not ( n77345 , n69587 );
not ( n77346 , n77345 );
not ( n77347 , n70308 );
or ( n77348 , n77346 , n77347 );
nand ( n77349 , n77348 , n77328 );
not ( n77350 , n70273 );
nand ( n77351 , n77350 , n69519 );
xor ( n77352 , n77349 , n77351 );
not ( n77353 , n69706 );
nand ( n77354 , n77353 , n77268 );
nand ( n77355 , n77270 , n77354 );
not ( n77356 , n72534 );
nand ( n77357 , n77356 , n69685 );
xor ( n77358 , n77355 , n77357 );
not ( n77359 , n69685 );
nand ( n77360 , n77359 , n72534 );
nand ( n77361 , n77357 , n77360 );
xor ( n77362 , n77361 , n77340 );
nand ( n77363 , n77344 , n77352 , n77358 , n77362 );
nor ( n77364 , n77338 , n77363 );
not ( n77365 , n69655 );
nand ( n77366 , n77365 , n71074 );
nand ( n77367 , n77314 , n77366 );
and ( n77368 , n77367 , n77243 );
not ( n77369 , n77367 );
not ( n77370 , n77243 );
and ( n77371 , n77369 , n77370 );
nor ( n77372 , n77368 , n77371 );
not ( n77373 , n69896 );
nand ( n77374 , n77373 , n72475 );
nand ( n77375 , n77336 , n77374 );
not ( n77376 , n72485 );
nand ( n77377 , n77376 , n69871 );
xor ( n77378 , n77375 , n77377 );
not ( n77379 , n70273 );
not ( n77380 , n69519 );
not ( n77381 , n77380 );
or ( n77382 , n77379 , n77381 );
nand ( n77383 , n77382 , n77351 );
not ( n77384 , n70253 );
nand ( n77385 , n77384 , n69531 );
xor ( n77386 , n77383 , n77385 );
not ( n77387 , n69435 );
not ( n77388 , n77387 );
not ( n77389 , n70477 );
or ( n77390 , n77388 , n77389 );
not ( n77391 , n70477 );
nand ( n77392 , n77391 , n69435 );
nand ( n77393 , n77390 , n77392 );
not ( n77394 , n70432 );
nand ( n77395 , n77394 , n69502 );
xor ( n77396 , n77393 , n77395 );
nand ( n77397 , n77372 , n77378 , n77386 , n77396 );
not ( n77398 , n70327 );
not ( n77399 , n69599 );
not ( n77400 , n77399 );
or ( n77401 , n77398 , n77400 );
not ( n77402 , n70327 );
nand ( n77403 , n77402 , n69599 );
nand ( n77404 , n77401 , n77403 );
xor ( n77405 , n77404 , n77325 );
not ( n77406 , n70238 );
not ( n77407 , n69613 );
not ( n77408 , n77407 );
or ( n77409 , n77406 , n77408 );
nand ( n77410 , n77409 , n77248 );
xor ( n77411 , n77410 , n77403 );
not ( n77412 , n69871 );
nand ( n77413 , n77412 , n72485 );
nand ( n77414 , n77377 , n77413 );
xor ( n77415 , n77414 , n77299 );
not ( n77416 , n69769 );
nand ( n77417 , n77416 , n72510 );
nand ( n77418 , n77260 , n77417 );
xor ( n77419 , n77418 , n77331 );
nand ( n77420 , n77405 , n77411 , n77415 , n77419 );
nor ( n77421 , n77397 , n77420 );
not ( n77422 , n69743 );
nand ( n77423 , n77422 , n73916 );
nand ( n77424 , n77273 , n77423 );
xor ( n77425 , n77424 , n77264 );
not ( n77426 , n69487 );
not ( n77427 , n77426 );
not ( n77428 , n70817 );
not ( n77429 , n77428 );
or ( n77430 , n77427 , n77429 );
not ( n77431 , n77428 );
nand ( n77432 , n77431 , n69487 );
nand ( n77433 , n77430 , n77432 );
not ( n77434 , n70420 );
nand ( n77435 , n77434 , n69471 );
xor ( n77436 , n77433 , n77435 );
not ( n77437 , n69470 );
not ( n77438 , n77437 );
not ( n77439 , n70388 );
or ( n77440 , n77438 , n77439 );
not ( n77441 , n70388 );
nand ( n77442 , n77441 , n69470 );
nand ( n77443 , n77440 , n77442 );
xor ( n77444 , n77443 , n77392 );
not ( n77445 , n69543 );
not ( n77446 , n77445 );
not ( n77447 , n70263 );
or ( n77448 , n77446 , n77447 );
not ( n77449 , n70263 );
nand ( n77450 , n77449 , n69543 );
nand ( n77451 , n77448 , n77450 );
not ( n77452 , n70378 );
nand ( n77453 , n77452 , n69553 );
xor ( n77454 , n77451 , n77453 );
nand ( n77455 , n77425 , n77436 , n77444 , n77454 );
not ( n77456 , n70253 );
not ( n77457 , n69531 );
not ( n77458 , n77457 );
or ( n77459 , n77456 , n77458 );
nand ( n77460 , n77459 , n77385 );
xor ( n77461 , n77460 , n77450 );
not ( n77462 , n69502 );
not ( n77463 , n77462 );
not ( n77464 , n70432 );
or ( n77465 , n77463 , n77464 );
nand ( n77466 , n77465 , n77395 );
and ( n77467 , n77466 , n77432 );
not ( n77468 , n77466 );
not ( n77469 , n77432 );
and ( n77470 , n77468 , n77469 );
nor ( n77471 , n77467 , n77470 );
not ( n77472 , n69553 );
not ( n77473 , n77472 );
not ( n77474 , n70378 );
or ( n77475 , n77473 , n77474 );
nand ( n77476 , n77475 , n77453 );
xor ( n77477 , n77476 , n77442 );
xnor ( n77478 , n70073 , n70459 );
not ( n77479 , n69967 );
and ( n77480 , n70522 , n77479 );
not ( n77481 , n70522 );
and ( n77482 , n77481 , n69967 );
nor ( n77483 , n77480 , n77482 );
xnor ( n77484 , n70503 , n70053 );
nand ( n77485 , n77478 , n77483 , n77484 );
xor ( n77486 , n69471 , n69451 );
xor ( n77487 , n77486 , n70420 );
nor ( n77488 , n77485 , n77487 );
nand ( n77489 , n77461 , n77471 , n77477 , n77488 );
nor ( n77490 , n77455 , n77489 );
and ( n77491 , n77293 , n77364 , n77421 , n77490 );
not ( n77492 , n70188 );
nor ( n77493 , n77492 , n70863 , n70194 );
not ( n77494 , n77493 );
or ( n77495 , n77491 , n77494 );
nand ( n77496 , n77493 , n70151 );
nand ( n77497 , n77495 , n77496 );
not ( n77498 , n77497 );
or ( n77499 , n77241 , n77498 );
nor ( n77500 , n70560 , n70863 );
nand ( n77501 , n77500 , n77240 );
nor ( n77502 , n77491 , n77501 );
not ( n77503 , n71983 );
nand ( n77504 , n70202 , n70865 , n70139 );
and ( n77505 , n70873 , n77503 , n77504 );
nor ( n77506 , n77505 , n77496 );
nor ( n77507 , n77502 , n77506 );
nand ( n77508 , n77499 , n77507 );
nor ( n77509 , n77239 , n77508 );
and ( n77510 , n77225 , n77234 , n77509 );
not ( n77511 , n71122 );
nor ( n77512 , n71058 , n77511 );
not ( n77513 , n71092 );
nor ( n77514 , n71047 , n77513 );
nor ( n77515 , n77512 , n77514 );
not ( n77516 , n71074 );
nand ( n77517 , n77516 , n69660 );
not ( n77518 , n70225 );
nand ( n77519 , n77518 , n69977 );
and ( n77520 , n77517 , n77519 );
not ( n77521 , n71074 );
nor ( n77522 , n77521 , n69660 );
nor ( n77523 , n77520 , n77522 );
and ( n77524 , n77515 , n77523 );
not ( n77525 , n71092 );
nand ( n77526 , n77525 , n71047 );
or ( n77527 , n77512 , n77526 );
nand ( n77528 , n71058 , n77511 );
nand ( n77529 , n77527 , n77528 );
nor ( n77530 , n77524 , n77529 );
not ( n77531 , n71833 );
not ( n77532 , n72510 );
nor ( n77533 , n77531 , n77532 );
not ( n77534 , n72499 );
nor ( n77535 , n71852 , n77534 );
nor ( n77536 , n77533 , n77535 );
not ( n77537 , n72475 );
nor ( n77538 , n71869 , n77537 );
not ( n77539 , n72485 );
nor ( n77540 , n77539 , n71037 );
nor ( n77541 , n77538 , n77540 );
nand ( n77542 , n77536 , n77541 );
or ( n77543 , n77530 , n77542 );
not ( n77544 , n71869 );
not ( n77545 , n77537 );
or ( n77546 , n77544 , n77545 );
not ( n77547 , n72485 );
nand ( n77548 , n77547 , n71037 );
or ( n77549 , n77538 , n77548 );
nand ( n77550 , n77546 , n77549 );
and ( n77551 , n77550 , n77536 );
nand ( n77552 , n71852 , n77534 );
or ( n77553 , n77533 , n77552 );
nand ( n77554 , n77531 , n77532 );
nand ( n77555 , n77553 , n77554 );
nor ( n77556 , n77551 , n77555 );
nand ( n77557 , n77543 , n77556 );
not ( n77558 , n77557 );
not ( n77559 , n73914 );
not ( n77560 , n73902 );
not ( n77561 , n77560 );
or ( n77562 , n77559 , n77561 );
not ( n77563 , n73912 );
nand ( n77564 , n69947 , n77563 );
nand ( n77565 , n77562 , n77564 );
not ( n77566 , n77565 );
not ( n77567 , n73916 );
nor ( n77568 , n72463 , n77567 );
not ( n77569 , n72626 );
nor ( n77570 , n77569 , n72452 );
nor ( n77571 , n77568 , n77570 );
nand ( n77572 , n77566 , n77571 );
not ( n77573 , n72815 );
nor ( n77574 , n77573 , n71763 );
not ( n77575 , n72534 );
nor ( n77576 , n77575 , n76748 );
nor ( n77577 , n77574 , n77576 );
not ( n77578 , n72544 );
nor ( n77579 , n76781 , n77578 );
not ( n77580 , n72557 );
nor ( n77581 , n71814 , n77580 );
nor ( n77582 , n77579 , n77581 );
nand ( n77583 , n77577 , n77582 );
nor ( n77584 , n77572 , n77583 );
not ( n77585 , n77584 );
or ( n77586 , n77558 , n77585 );
not ( n77587 , n77572 );
nand ( n77588 , n76781 , n77578 );
nand ( n77589 , n71814 , n77580 );
and ( n77590 , n77588 , n77589 );
nor ( n77591 , n77590 , n77579 );
not ( n77592 , n77591 );
not ( n77593 , n77577 );
or ( n77594 , n77592 , n77593 );
not ( n77595 , n77574 );
not ( n77596 , n76748 );
nor ( n77597 , n77596 , n72534 );
and ( n77598 , n77595 , n77597 );
not ( n77599 , n71763 );
nor ( n77600 , n77599 , n72815 );
nor ( n77601 , n77598 , n77600 );
nand ( n77602 , n77594 , n77601 );
and ( n77603 , n77587 , n77602 );
not ( n77604 , n72463 );
not ( n77605 , n77604 );
not ( n77606 , n73916 );
and ( n77607 , n77605 , n77606 );
not ( n77608 , n77568 );
not ( n77609 , n72452 );
nor ( n77610 , n77609 , n72626 );
and ( n77611 , n77608 , n77610 );
nor ( n77612 , n77607 , n77611 );
or ( n77613 , n77612 , n77565 );
not ( n77614 , n73902 );
nor ( n77615 , n77614 , n73914 );
and ( n77616 , n77564 , n77615 );
nor ( n77617 , n69947 , n77563 );
nor ( n77618 , n77616 , n77617 );
nand ( n77619 , n77613 , n77618 );
nor ( n77620 , n77603 , n77619 );
nand ( n77621 , n77586 , n77620 );
not ( n77622 , n76395 );
nand ( n77623 , n77622 , n70238 );
not ( n77624 , n69981 );
nand ( n77625 , n77624 , n70327 );
nand ( n77626 , n77623 , n77625 );
not ( n77627 , n70098 );
nand ( n77628 , n77627 , n70296 );
not ( n77629 , n69990 );
nand ( n77630 , n77629 , n70308 );
nand ( n77631 , n77628 , n77630 );
nor ( n77632 , n77626 , n77631 );
not ( n77633 , n70273 );
nor ( n77634 , n77633 , n76513 );
not ( n77635 , n70253 );
nor ( n77636 , n77635 , n70013 );
nor ( n77637 , n77634 , n77636 );
not ( n77638 , n77637 );
not ( n77639 , n70378 );
not ( n77640 , n70082 );
not ( n77641 , n77640 );
or ( n77642 , n77639 , n77641 );
not ( n77643 , n70263 );
nor ( n77644 , n77643 , n70007 );
not ( n77645 , n77644 );
nand ( n77646 , n77642 , n77645 );
nor ( n77647 , n77638 , n77646 );
not ( n77648 , n70388 );
nor ( n77649 , n77648 , n70090 );
not ( n77650 , n70477 );
nor ( n77651 , n77650 , n70031 );
nor ( n77652 , n77649 , n77651 );
not ( n77653 , n70432 );
nor ( n77654 , n70024 , n77653 );
not ( n77655 , n72302 );
nor ( n77656 , n77655 , n70038 );
nor ( n77657 , n77654 , n77656 );
not ( n77658 , n70040 );
nand ( n77659 , n77658 , n70420 );
not ( n77660 , n70522 );
nor ( n77661 , n77660 , n69967 );
not ( n77662 , n70053 );
and ( n77663 , n77662 , n70503 );
or ( n77664 , n77661 , n77663 );
or ( n77665 , n77662 , n70503 );
nand ( n77666 , n77664 , n77665 );
not ( n77667 , n70073 );
nand ( n77668 , n77667 , n70459 );
nand ( n77669 , n77659 , n77666 , n77668 );
not ( n77670 , n70073 );
nor ( n77671 , n77670 , n70459 );
nand ( n77672 , n77659 , n77671 );
not ( n77673 , n70420 );
nand ( n77674 , n77673 , n70040 );
nand ( n77675 , n77669 , n77672 , n77674 );
nand ( n77676 , n77652 , n77657 , n77675 );
not ( n77677 , n72302 );
nand ( n77678 , n77677 , n70038 );
or ( n77679 , n77654 , n77678 );
nand ( n77680 , n70024 , n77653 );
nand ( n77681 , n77679 , n77680 );
nand ( n77682 , n77652 , n77681 );
not ( n77683 , n77649 );
not ( n77684 , n70031 );
nor ( n77685 , n77684 , n70477 );
and ( n77686 , n77683 , n77685 );
not ( n77687 , n70090 );
nor ( n77688 , n77687 , n70388 );
nor ( n77689 , n77686 , n77688 );
nand ( n77690 , n77676 , n77682 , n77689 );
nand ( n77691 , n77632 , n77647 , n77690 );
not ( n77692 , n77637 );
not ( n77693 , n70378 );
nand ( n77694 , n77693 , n70082 );
or ( n77695 , n77644 , n77694 );
not ( n77696 , n70007 );
or ( n77697 , n77696 , n70263 );
nand ( n77698 , n77695 , n77697 );
not ( n77699 , n77698 );
or ( n77700 , n77692 , n77699 );
not ( n77701 , n77634 );
not ( n77702 , n70013 );
nor ( n77703 , n77702 , n70253 );
and ( n77704 , n77701 , n77703 );
not ( n77705 , n76513 );
nor ( n77706 , n77705 , n70273 );
nor ( n77707 , n77704 , n77706 );
nand ( n77708 , n77700 , n77707 );
nand ( n77709 , n77708 , n77632 );
not ( n77710 , n77628 );
not ( n77711 , n70308 );
nand ( n77712 , n77711 , n69990 );
or ( n77713 , n77710 , n77712 );
not ( n77714 , n70296 );
nand ( n77715 , n77714 , n70098 );
nand ( n77716 , n77713 , n77715 );
not ( n77717 , n77626 );
and ( n77718 , n77716 , n77717 );
not ( n77719 , n77623 );
not ( n77720 , n70327 );
nand ( n77721 , n77720 , n69981 );
or ( n77722 , n77719 , n77721 );
not ( n77723 , n70238 );
nand ( n77724 , n77723 , n76395 );
nand ( n77725 , n77722 , n77724 );
nor ( n77726 , n77718 , n77725 );
nand ( n77727 , n77691 , n77709 , n77726 );
not ( n77728 , n70225 );
nor ( n77729 , n77728 , n69977 );
nor ( n77730 , n77522 , n77729 );
nand ( n77731 , n77515 , n77730 );
nor ( n77732 , n77542 , n77731 );
not ( n77733 , n77583 );
and ( n77734 , n77587 , n77727 , n77732 , n77733 );
nor ( n77735 , n77621 , n77734 );
or ( n77736 , n77735 , n70873 );
not ( n77737 , n77504 );
nand ( n77738 , n77491 , n77737 );
nand ( n77739 , n77736 , n77738 );
not ( n77740 , n77739 );
nand ( n77741 , n77735 , n71983 );
nand ( n77742 , n77740 , n77741 );
nand ( n77743 , n77742 , n77493 );
nand ( n77744 , n77742 , n77500 );
and ( n77745 , n77229 , n77737 );
not ( n77746 , n77223 );
and ( n77747 , n77746 , n77240 );
nor ( n77748 , n77745 , n77747 );
and ( n77749 , n77510 , n77743 , n77744 , n77748 );
or ( n77750 , n76991 , n77749 );
nand ( n77751 , n77510 , n77743 , n77744 );
not ( n77752 , n77240 );
not ( n77753 , n77229 );
or ( n77754 , n77752 , n77753 );
or ( n77755 , n77223 , n77504 );
nand ( n77756 , n77754 , n77755 );
nor ( n77757 , n77751 , n77756 );
or ( n77758 , n77757 , n76990 );
not ( n77759 , n75275 );
nor ( n77760 , n70141 , n70208 , n77759 );
not ( n77761 , n77760 );
nand ( n77762 , n70147 , n70860 );
nand ( n77763 , n77761 , n77762 , n70151 );
nand ( n77764 , n77750 , n77758 , n77763 );
buf ( n77765 , n77764 );
buf ( n77766 , 1'b0 );
not ( n77767 , n68635 );
not ( n77768 , n77767 );
buf ( n77769 , n77768 );
buf ( n77770 , n68634 );
buf ( n77771 , n71724 );
buf ( n77772 , 1'b0 );
not ( n77773 , n77767 );
buf ( n77774 , n77773 );
buf ( n77775 , n68634 );
nand ( n77776 , n70188 , n70194 );
and ( n77777 , n70136 , n77776 );
nor ( n77778 , n77777 , n70147 );
not ( n77779 , n70222 );
or ( n77780 , n77778 , n77779 );
nand ( n77781 , n77780 , n70860 );
buf ( n77782 , n77781 );
endmodule
